// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"

// DATE "01/25/2021 23:31:52"

// 
// Device: Altera 5CSXFC6D6F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module soc_system (
	clk_clk,
	clk_100m_clk,
	d_out_in,
	d_out_out,
	d_out_oe,
	hps_io_hps_io_emac1_inst_TX_CLK,
	hps_io_hps_io_emac1_inst_TXD0,
	hps_io_hps_io_emac1_inst_TXD1,
	hps_io_hps_io_emac1_inst_TXD2,
	hps_io_hps_io_emac1_inst_TXD3,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_MDIO,
	hps_io_hps_io_emac1_inst_MDC,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_emac1_inst_TX_CTL,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_qspi_inst_IO0,
	hps_io_hps_io_qspi_inst_IO1,
	hps_io_hps_io_qspi_inst_IO2,
	hps_io_hps_io_qspi_inst_IO3,
	hps_io_hps_io_qspi_inst_SS0,
	hps_io_hps_io_qspi_inst_CLK,
	hps_io_hps_io_sdio_inst_CMD,
	hps_io_hps_io_sdio_inst_D0,
	hps_io_hps_io_sdio_inst_D1,
	hps_io_hps_io_sdio_inst_CLK,
	hps_io_hps_io_sdio_inst_D2,
	hps_io_hps_io_sdio_inst_D3,
	hps_io_hps_io_usb1_inst_D0,
	hps_io_hps_io_usb1_inst_D1,
	hps_io_hps_io_usb1_inst_D2,
	hps_io_hps_io_usb1_inst_D3,
	hps_io_hps_io_usb1_inst_D4,
	hps_io_hps_io_usb1_inst_D5,
	hps_io_hps_io_usb1_inst_D6,
	hps_io_hps_io_usb1_inst_D7,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_STP,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	hps_io_hps_io_spim0_inst_CLK,
	hps_io_hps_io_spim0_inst_MOSI,
	hps_io_hps_io_spim0_inst_MISO,
	hps_io_hps_io_spim0_inst_SS0,
	hps_io_hps_io_spim1_inst_CLK,
	hps_io_hps_io_spim1_inst_MOSI,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_spim1_inst_SS0,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_uart0_inst_TX,
	hps_io_hps_io_gpio_inst_GPIO09,
	hps_io_hps_io_gpio_inst_GPIO40,
	hps_io_hps_io_gpio_inst_GPIO48,
	hps_io_hps_io_gpio_inst_GPIO61,
	hps_io_hps_io_gpio_inst_GPIO62,
	hps_io_hps_io_gpio_inst_LOANIO00,
	hps_io_hps_io_gpio_inst_LOANIO41,
	hps_io_hps_io_gpio_inst_LOANIO51,
	hps_io_hps_io_gpio_inst_LOANIO52,
	hps_io_hps_io_gpio_inst_LOANIO53,
	hps_io_hps_io_gpio_inst_LOANIO54,
	hps_io_hps_io_gpio_inst_LOANIO55,
	hps_io_hps_io_gpio_inst_LOANIO56,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	ram_clk_clk,
	ram_mm_address,
	ram_mm_chipselect,
	ram_mm_clken,
	ram_mm_write,
	ram_mm_readdata,
	ram_mm_writedata,
	ram_mm_byteenable,
	ram_reset_reset,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	clk_clk;
output 	clk_100m_clk;
output 	[66:0] d_out_in;
input 	[66:0] d_out_out;
input 	[66:0] d_out_oe;
output 	hps_io_hps_io_emac1_inst_TX_CLK;
output 	hps_io_hps_io_emac1_inst_TXD0;
output 	hps_io_hps_io_emac1_inst_TXD1;
output 	hps_io_hps_io_emac1_inst_TXD2;
output 	hps_io_hps_io_emac1_inst_TXD3;
input 	hps_io_hps_io_emac1_inst_RXD0;
inout 	hps_io_hps_io_emac1_inst_MDIO;
output 	hps_io_hps_io_emac1_inst_MDC;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
output 	hps_io_hps_io_emac1_inst_TX_CTL;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
inout 	hps_io_hps_io_qspi_inst_IO0;
inout 	hps_io_hps_io_qspi_inst_IO1;
inout 	hps_io_hps_io_qspi_inst_IO2;
inout 	hps_io_hps_io_qspi_inst_IO3;
output 	hps_io_hps_io_qspi_inst_SS0;
output 	hps_io_hps_io_qspi_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_CMD;
inout 	hps_io_hps_io_sdio_inst_D0;
inout 	hps_io_hps_io_sdio_inst_D1;
output 	hps_io_hps_io_sdio_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_D2;
inout 	hps_io_hps_io_sdio_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D0;
inout 	hps_io_hps_io_usb1_inst_D1;
inout 	hps_io_hps_io_usb1_inst_D2;
inout 	hps_io_hps_io_usb1_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D4;
inout 	hps_io_hps_io_usb1_inst_D5;
inout 	hps_io_hps_io_usb1_inst_D6;
inout 	hps_io_hps_io_usb1_inst_D7;
input 	hps_io_hps_io_usb1_inst_CLK;
output 	hps_io_hps_io_usb1_inst_STP;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
output 	hps_io_hps_io_spim0_inst_CLK;
output 	hps_io_hps_io_spim0_inst_MOSI;
input 	hps_io_hps_io_spim0_inst_MISO;
output 	hps_io_hps_io_spim0_inst_SS0;
output 	hps_io_hps_io_spim1_inst_CLK;
output 	hps_io_hps_io_spim1_inst_MOSI;
input 	hps_io_hps_io_spim1_inst_MISO;
output 	hps_io_hps_io_spim1_inst_SS0;
input 	hps_io_hps_io_uart0_inst_RX;
output 	hps_io_hps_io_uart0_inst_TX;
inout 	hps_io_hps_io_gpio_inst_GPIO09;
inout 	hps_io_hps_io_gpio_inst_GPIO40;
inout 	hps_io_hps_io_gpio_inst_GPIO48;
inout 	hps_io_hps_io_gpio_inst_GPIO61;
inout 	hps_io_hps_io_gpio_inst_GPIO62;
inout 	hps_io_hps_io_gpio_inst_LOANIO00;
inout 	hps_io_hps_io_gpio_inst_LOANIO41;
inout 	hps_io_hps_io_gpio_inst_LOANIO51;
inout 	hps_io_hps_io_gpio_inst_LOANIO52;
inout 	hps_io_hps_io_gpio_inst_LOANIO53;
inout 	hps_io_hps_io_gpio_inst_LOANIO54;
inout 	hps_io_hps_io_gpio_inst_LOANIO55;
inout 	hps_io_hps_io_gpio_inst_LOANIO56;
output 	[14:0] memory_mem_a;
output 	[2:0] memory_mem_ba;
output 	memory_mem_ck;
output 	memory_mem_ck_n;
output 	memory_mem_cke;
output 	memory_mem_cs_n;
output 	memory_mem_ras_n;
output 	memory_mem_cas_n;
output 	memory_mem_we_n;
output 	memory_mem_reset_n;
inout 	[31:0] memory_mem_dq;
inout 	[3:0] memory_mem_dqs;
inout 	[3:0] memory_mem_dqs_n;
output 	memory_mem_odt;
output 	[3:0] memory_mem_dm;
input 	memory_oct_rzqin;
input 	ram_clk_clk;
input 	[12:0] ram_mm_address;
input 	ram_mm_chipselect;
input 	ram_mm_clken;
input 	ram_mm_write;
output 	[31:0] ram_mm_readdata;
input 	[31:0] ram_mm_writedata;
input 	[3:0] ram_mm_byteenable;
input 	ram_reset_reset;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0|fpga_interfaces|h2f_loan_in[0] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[1] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[2] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[3] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[4] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[5] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[6] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[7] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[8] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[9] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[10] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[11] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[12] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[13] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[14] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[15] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[16] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[17] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[18] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[19] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[20] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[21] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[22] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[23] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[24] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[25] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[26] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[27] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[28] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[29] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[30] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[31] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[32] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[33] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[34] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[35] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[36] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[37] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[38] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[39] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[40] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[41] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[42] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[43] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[44] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[45] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[46] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[47] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[48] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[49] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[50] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[51] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[52] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[53] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[54] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[55] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[56] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[57] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[58] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[59] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[60] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[61] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[62] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[63] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[64] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[65] ;
wire \hps_0|fpga_interfaces|h2f_loan_in[66] ;
wire \hps_0|fpga_interfaces|h2f_rst_n[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_BREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_RREADY[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WLAST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WVALID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[12] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[13] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARADDR[14] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARID[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[12] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[13] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWADDR[14] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWID[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[3] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[4] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[5] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[6] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[7] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[8] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[9] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[10] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[11] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[12] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[13] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[14] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[15] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[16] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[17] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[18] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[19] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[20] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[21] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[22] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[23] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[24] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[25] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[26] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[27] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[28] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[29] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[30] ;
wire \hps_0|fpga_interfaces|h2f_lw_WDATA[31] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ;
wire \hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ;
wire \pll_0|altera_pll_i|outclk_wire[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[16] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[17] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[18] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[19] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_b[31] ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~2_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~3_combout ;
wire \mm_interconnect_0|cmd_mux|sink1_ready~combout ;
wire \mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ;
wire \mm_interconnect_0|rsp_demux|src0_valid~combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent|uncompressor|source_endofpacket~combout ;
wire \mm_interconnect_0|rsp_demux|src1_valid~0_combout ;
wire \mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][88]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][89]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][90]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][91]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[0]~0_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[1]~1_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[2]~2_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[3]~3_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[4]~4_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[5]~5_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[6]~6_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[7]~7_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[8]~8_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[9]~9_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[10]~10_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[11]~11_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[12]~12_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[13]~13_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[14]~14_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[15]~15_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[16]~16_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[17]~17_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[18]~18_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[19]~19_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[20]~20_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[21]~21_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[22]~22_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[23]~23_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[24]~24_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[25]~25_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[26]~26_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[27]~27_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[28]~28_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[29]~29_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[30]~30_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[31]~31_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent|m0_write~1_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[10]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[11]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[12]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[13]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[14]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~7_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~8_combout ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;
wire \hps_0|hps_io|border|intermediate[0] ;
wire \hps_0|hps_io|border|intermediate[1] ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;
wire \hps_0|hps_io|border|emac1_inst~emac_phy_txd ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;
wire \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;
wire \hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ;
wire \hps_0|hps_io|border|intermediate[2] ;
wire \hps_0|hps_io|border|intermediate[4] ;
wire \hps_0|hps_io|border|intermediate[6] ;
wire \hps_0|hps_io|border|intermediate[8] ;
wire \hps_0|hps_io|border|intermediate[3] ;
wire \hps_0|hps_io|border|intermediate[5] ;
wire \hps_0|hps_io|border|intermediate[7] ;
wire \hps_0|hps_io|border|intermediate[9] ;
wire \hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;
wire \hps_0|hps_io|border|sdio_inst~sdmmc_cclk ;
wire \hps_0|hps_io|border|intermediate[10] ;
wire \hps_0|hps_io|border|intermediate[11] ;
wire \hps_0|hps_io|border|intermediate[12] ;
wire \hps_0|hps_io|border|intermediate[14] ;
wire \hps_0|hps_io|border|intermediate[16] ;
wire \hps_0|hps_io|border|intermediate[18] ;
wire \hps_0|hps_io|border|intermediate[13] ;
wire \hps_0|hps_io|border|intermediate[15] ;
wire \hps_0|hps_io|border|intermediate[17] ;
wire \hps_0|hps_io|border|intermediate[19] ;
wire \hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ;
wire \hps_0|hps_io|border|intermediate[20] ;
wire \hps_0|hps_io|border|intermediate[22] ;
wire \hps_0|hps_io|border|intermediate[24] ;
wire \hps_0|hps_io|border|intermediate[26] ;
wire \hps_0|hps_io|border|intermediate[28] ;
wire \hps_0|hps_io|border|intermediate[30] ;
wire \hps_0|hps_io|border|intermediate[32] ;
wire \hps_0|hps_io|border|intermediate[34] ;
wire \hps_0|hps_io|border|intermediate[21] ;
wire \hps_0|hps_io|border|intermediate[23] ;
wire \hps_0|hps_io|border|intermediate[25] ;
wire \hps_0|hps_io|border|intermediate[27] ;
wire \hps_0|hps_io|border|intermediate[29] ;
wire \hps_0|hps_io|border|intermediate[31] ;
wire \hps_0|hps_io|border|intermediate[33] ;
wire \hps_0|hps_io|border|intermediate[35] ;
wire \hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SCLK ;
wire \hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SS_0_N ;
wire \hps_0|hps_io|border|intermediate[36] ;
wire \hps_0|hps_io|border|intermediate[37] ;
wire \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;
wire \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;
wire \hps_0|hps_io|border|intermediate[38] ;
wire \hps_0|hps_io|border|intermediate[39] ;
wire \hps_0|hps_io|border|uart0_inst~uart_txd ;
wire \hps_0|hps_io|border|intermediate[50] ;
wire \hps_0|hps_io|border|intermediate[40] ;
wire \hps_0|hps_io|border|intermediate[51] ;
wire \hps_0|hps_io|border|intermediate[41] ;
wire \hps_0|hps_io|border|intermediate[42] ;
wire \hps_0|hps_io|border|intermediate[52] ;
wire \hps_0|hps_io|border|intermediate[44] ;
wire \hps_0|hps_io|border|intermediate[54] ;
wire \hps_0|hps_io|border|intermediate[56] ;
wire \hps_0|hps_io|border|intermediate[58] ;
wire \hps_0|hps_io|border|intermediate[60] ;
wire \hps_0|hps_io|border|intermediate[62] ;
wire \hps_0|hps_io|border|intermediate[64] ;
wire \hps_0|hps_io|border|intermediate[43] ;
wire \hps_0|hps_io|border|intermediate[53] ;
wire \hps_0|hps_io|border|intermediate[45] ;
wire \hps_0|hps_io|border|intermediate[55] ;
wire \hps_0|hps_io|border|intermediate[57] ;
wire \hps_0|hps_io|border|intermediate[59] ;
wire \hps_0|hps_io|border|intermediate[61] ;
wire \hps_0|hps_io|border|intermediate[63] ;
wire \hps_0|hps_io|border|intermediate[65] ;
wire \hps_0|hps_io|border|intermediate[46] ;
wire \hps_0|hps_io|border|intermediate[48] ;
wire \hps_0|hps_io|border|intermediate[47] ;
wire \hps_0|hps_io|border|intermediate[49] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \ram_reset_reset~input_o ;
wire \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~input_o ;
wire \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD0~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD1~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD2~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD3~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CLK~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CTL~input_o ;
wire \hps_io_hps_io_spim0_inst_MISO~input_o ;
wire \hps_io_hps_io_spim1_inst_MISO~input_o ;
wire \hps_io_hps_io_uart0_inst_RX~input_o ;
wire \hps_io_hps_io_usb1_inst_CLK~input_o ;
wire \hps_io_hps_io_usb1_inst_DIR~input_o ;
wire \hps_io_hps_io_usb1_inst_NXT~input_o ;
wire \memory_oct_rzqin~input_o ;
wire \d_out_oe[0]~input_o ;
wire \d_out_oe[1]~input_o ;
wire \d_out_oe[2]~input_o ;
wire \d_out_oe[3]~input_o ;
wire \d_out_oe[4]~input_o ;
wire \d_out_oe[5]~input_o ;
wire \d_out_oe[6]~input_o ;
wire \d_out_oe[7]~input_o ;
wire \d_out_oe[8]~input_o ;
wire \d_out_oe[9]~input_o ;
wire \d_out_oe[10]~input_o ;
wire \d_out_oe[11]~input_o ;
wire \d_out_oe[12]~input_o ;
wire \d_out_oe[13]~input_o ;
wire \d_out_oe[14]~input_o ;
wire \d_out_oe[15]~input_o ;
wire \d_out_oe[16]~input_o ;
wire \d_out_oe[17]~input_o ;
wire \d_out_oe[18]~input_o ;
wire \d_out_oe[19]~input_o ;
wire \d_out_oe[20]~input_o ;
wire \d_out_oe[21]~input_o ;
wire \d_out_oe[22]~input_o ;
wire \d_out_oe[23]~input_o ;
wire \d_out_oe[24]~input_o ;
wire \d_out_oe[25]~input_o ;
wire \d_out_oe[26]~input_o ;
wire \d_out_oe[27]~input_o ;
wire \d_out_oe[28]~input_o ;
wire \d_out_oe[29]~input_o ;
wire \d_out_oe[30]~input_o ;
wire \d_out_oe[31]~input_o ;
wire \d_out_oe[32]~input_o ;
wire \d_out_oe[33]~input_o ;
wire \d_out_oe[34]~input_o ;
wire \d_out_oe[35]~input_o ;
wire \d_out_oe[36]~input_o ;
wire \d_out_oe[37]~input_o ;
wire \d_out_oe[38]~input_o ;
wire \d_out_oe[39]~input_o ;
wire \d_out_oe[40]~input_o ;
wire \d_out_oe[41]~input_o ;
wire \d_out_oe[42]~input_o ;
wire \d_out_oe[43]~input_o ;
wire \d_out_oe[44]~input_o ;
wire \d_out_oe[45]~input_o ;
wire \d_out_oe[46]~input_o ;
wire \d_out_oe[47]~input_o ;
wire \d_out_oe[48]~input_o ;
wire \d_out_oe[49]~input_o ;
wire \d_out_oe[50]~input_o ;
wire \d_out_oe[51]~input_o ;
wire \d_out_oe[52]~input_o ;
wire \d_out_oe[53]~input_o ;
wire \d_out_oe[54]~input_o ;
wire \d_out_oe[55]~input_o ;
wire \d_out_oe[56]~input_o ;
wire \d_out_oe[57]~input_o ;
wire \d_out_oe[58]~input_o ;
wire \d_out_oe[59]~input_o ;
wire \d_out_oe[60]~input_o ;
wire \d_out_oe[61]~input_o ;
wire \d_out_oe[62]~input_o ;
wire \d_out_oe[63]~input_o ;
wire \d_out_oe[64]~input_o ;
wire \d_out_oe[65]~input_o ;
wire \d_out_oe[66]~input_o ;
wire \d_out_out[0]~input_o ;
wire \d_out_out[1]~input_o ;
wire \d_out_out[2]~input_o ;
wire \d_out_out[3]~input_o ;
wire \d_out_out[4]~input_o ;
wire \d_out_out[5]~input_o ;
wire \d_out_out[6]~input_o ;
wire \d_out_out[7]~input_o ;
wire \d_out_out[8]~input_o ;
wire \d_out_out[9]~input_o ;
wire \d_out_out[10]~input_o ;
wire \d_out_out[11]~input_o ;
wire \d_out_out[12]~input_o ;
wire \d_out_out[13]~input_o ;
wire \d_out_out[14]~input_o ;
wire \d_out_out[15]~input_o ;
wire \d_out_out[16]~input_o ;
wire \d_out_out[17]~input_o ;
wire \d_out_out[18]~input_o ;
wire \d_out_out[19]~input_o ;
wire \d_out_out[20]~input_o ;
wire \d_out_out[21]~input_o ;
wire \d_out_out[22]~input_o ;
wire \d_out_out[23]~input_o ;
wire \d_out_out[24]~input_o ;
wire \d_out_out[25]~input_o ;
wire \d_out_out[26]~input_o ;
wire \d_out_out[27]~input_o ;
wire \d_out_out[28]~input_o ;
wire \d_out_out[29]~input_o ;
wire \d_out_out[30]~input_o ;
wire \d_out_out[31]~input_o ;
wire \d_out_out[32]~input_o ;
wire \d_out_out[33]~input_o ;
wire \d_out_out[34]~input_o ;
wire \d_out_out[35]~input_o ;
wire \d_out_out[36]~input_o ;
wire \d_out_out[37]~input_o ;
wire \d_out_out[38]~input_o ;
wire \d_out_out[39]~input_o ;
wire \d_out_out[40]~input_o ;
wire \d_out_out[41]~input_o ;
wire \d_out_out[42]~input_o ;
wire \d_out_out[43]~input_o ;
wire \d_out_out[44]~input_o ;
wire \d_out_out[45]~input_o ;
wire \d_out_out[46]~input_o ;
wire \d_out_out[47]~input_o ;
wire \d_out_out[48]~input_o ;
wire \d_out_out[49]~input_o ;
wire \d_out_out[50]~input_o ;
wire \d_out_out[51]~input_o ;
wire \d_out_out[52]~input_o ;
wire \d_out_out[53]~input_o ;
wire \d_out_out[54]~input_o ;
wire \d_out_out[55]~input_o ;
wire \d_out_out[56]~input_o ;
wire \d_out_out[57]~input_o ;
wire \d_out_out[58]~input_o ;
wire \d_out_out[59]~input_o ;
wire \d_out_out[60]~input_o ;
wire \d_out_out[61]~input_o ;
wire \d_out_out[62]~input_o ;
wire \d_out_out[63]~input_o ;
wire \d_out_out[64]~input_o ;
wire \d_out_out[65]~input_o ;
wire \d_out_out[66]~input_o ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \ram_mm_chipselect~input_o ;
wire \ram_mm_write~input_o ;
wire \ram_clk_clk~input_o ;
wire \ram_mm_clken~input_o ;
wire \ram_mm_writedata[0]~input_o ;
wire \ram_mm_address[0]~input_o ;
wire \ram_mm_address[1]~input_o ;
wire \ram_mm_address[2]~input_o ;
wire \ram_mm_address[3]~input_o ;
wire \ram_mm_address[4]~input_o ;
wire \ram_mm_address[5]~input_o ;
wire \ram_mm_address[6]~input_o ;
wire \ram_mm_address[7]~input_o ;
wire \ram_mm_address[8]~input_o ;
wire \ram_mm_address[9]~input_o ;
wire \ram_mm_address[10]~input_o ;
wire \ram_mm_address[11]~input_o ;
wire \ram_mm_address[12]~input_o ;
wire \ram_mm_byteenable[0]~input_o ;
wire \ram_mm_writedata[1]~input_o ;
wire \ram_mm_writedata[2]~input_o ;
wire \ram_mm_writedata[3]~input_o ;
wire \ram_mm_writedata[4]~input_o ;
wire \ram_mm_writedata[5]~input_o ;
wire \ram_mm_writedata[6]~input_o ;
wire \ram_mm_writedata[7]~input_o ;
wire \ram_mm_writedata[8]~input_o ;
wire \ram_mm_byteenable[1]~input_o ;
wire \ram_mm_writedata[9]~input_o ;
wire \ram_mm_writedata[10]~input_o ;
wire \ram_mm_writedata[11]~input_o ;
wire \ram_mm_writedata[12]~input_o ;
wire \ram_mm_writedata[13]~input_o ;
wire \ram_mm_writedata[14]~input_o ;
wire \ram_mm_writedata[15]~input_o ;
wire \ram_mm_writedata[16]~input_o ;
wire \ram_mm_byteenable[2]~input_o ;
wire \ram_mm_writedata[17]~input_o ;
wire \ram_mm_writedata[18]~input_o ;
wire \ram_mm_writedata[19]~input_o ;
wire \ram_mm_writedata[20]~input_o ;
wire \ram_mm_writedata[21]~input_o ;
wire \ram_mm_writedata[22]~input_o ;
wire \ram_mm_writedata[23]~input_o ;
wire \ram_mm_writedata[24]~input_o ;
wire \ram_mm_byteenable[3]~input_o ;
wire \ram_mm_writedata[25]~input_o ;
wire \ram_mm_writedata[26]~input_o ;
wire \ram_mm_writedata[27]~input_o ;
wire \ram_mm_writedata[28]~input_o ;
wire \ram_mm_writedata[29]~input_o ;
wire \ram_mm_writedata[30]~input_o ;
wire \ram_mm_writedata[31]~input_o ;


soc_system_altera_reset_controller_1 rst_controller_001(
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

soc_system_altera_reset_controller rst_controller(
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.reset_reset_n(\reset_reset_n~input_o ));

soc_system_soc_system_hps_0 hps_0(
	.h2f_loan_in_0(\hps_0|fpga_interfaces|h2f_loan_in[0] ),
	.h2f_loan_in_1(\hps_0|fpga_interfaces|h2f_loan_in[1] ),
	.h2f_loan_in_2(\hps_0|fpga_interfaces|h2f_loan_in[2] ),
	.h2f_loan_in_3(\hps_0|fpga_interfaces|h2f_loan_in[3] ),
	.h2f_loan_in_4(\hps_0|fpga_interfaces|h2f_loan_in[4] ),
	.h2f_loan_in_5(\hps_0|fpga_interfaces|h2f_loan_in[5] ),
	.h2f_loan_in_6(\hps_0|fpga_interfaces|h2f_loan_in[6] ),
	.h2f_loan_in_7(\hps_0|fpga_interfaces|h2f_loan_in[7] ),
	.h2f_loan_in_8(\hps_0|fpga_interfaces|h2f_loan_in[8] ),
	.h2f_loan_in_9(\hps_0|fpga_interfaces|h2f_loan_in[9] ),
	.h2f_loan_in_10(\hps_0|fpga_interfaces|h2f_loan_in[10] ),
	.h2f_loan_in_11(\hps_0|fpga_interfaces|h2f_loan_in[11] ),
	.h2f_loan_in_12(\hps_0|fpga_interfaces|h2f_loan_in[12] ),
	.h2f_loan_in_13(\hps_0|fpga_interfaces|h2f_loan_in[13] ),
	.h2f_loan_in_14(\hps_0|fpga_interfaces|h2f_loan_in[14] ),
	.h2f_loan_in_15(\hps_0|fpga_interfaces|h2f_loan_in[15] ),
	.h2f_loan_in_16(\hps_0|fpga_interfaces|h2f_loan_in[16] ),
	.h2f_loan_in_17(\hps_0|fpga_interfaces|h2f_loan_in[17] ),
	.h2f_loan_in_18(\hps_0|fpga_interfaces|h2f_loan_in[18] ),
	.h2f_loan_in_19(\hps_0|fpga_interfaces|h2f_loan_in[19] ),
	.h2f_loan_in_20(\hps_0|fpga_interfaces|h2f_loan_in[20] ),
	.h2f_loan_in_21(\hps_0|fpga_interfaces|h2f_loan_in[21] ),
	.h2f_loan_in_22(\hps_0|fpga_interfaces|h2f_loan_in[22] ),
	.h2f_loan_in_23(\hps_0|fpga_interfaces|h2f_loan_in[23] ),
	.h2f_loan_in_24(\hps_0|fpga_interfaces|h2f_loan_in[24] ),
	.h2f_loan_in_25(\hps_0|fpga_interfaces|h2f_loan_in[25] ),
	.h2f_loan_in_26(\hps_0|fpga_interfaces|h2f_loan_in[26] ),
	.h2f_loan_in_27(\hps_0|fpga_interfaces|h2f_loan_in[27] ),
	.h2f_loan_in_28(\hps_0|fpga_interfaces|h2f_loan_in[28] ),
	.h2f_loan_in_29(\hps_0|fpga_interfaces|h2f_loan_in[29] ),
	.h2f_loan_in_30(\hps_0|fpga_interfaces|h2f_loan_in[30] ),
	.h2f_loan_in_31(\hps_0|fpga_interfaces|h2f_loan_in[31] ),
	.h2f_loan_in_32(\hps_0|fpga_interfaces|h2f_loan_in[32] ),
	.h2f_loan_in_33(\hps_0|fpga_interfaces|h2f_loan_in[33] ),
	.h2f_loan_in_34(\hps_0|fpga_interfaces|h2f_loan_in[34] ),
	.h2f_loan_in_35(\hps_0|fpga_interfaces|h2f_loan_in[35] ),
	.h2f_loan_in_36(\hps_0|fpga_interfaces|h2f_loan_in[36] ),
	.h2f_loan_in_37(\hps_0|fpga_interfaces|h2f_loan_in[37] ),
	.h2f_loan_in_38(\hps_0|fpga_interfaces|h2f_loan_in[38] ),
	.h2f_loan_in_39(\hps_0|fpga_interfaces|h2f_loan_in[39] ),
	.h2f_loan_in_40(\hps_0|fpga_interfaces|h2f_loan_in[40] ),
	.h2f_loan_in_41(\hps_0|fpga_interfaces|h2f_loan_in[41] ),
	.h2f_loan_in_42(\hps_0|fpga_interfaces|h2f_loan_in[42] ),
	.h2f_loan_in_43(\hps_0|fpga_interfaces|h2f_loan_in[43] ),
	.h2f_loan_in_44(\hps_0|fpga_interfaces|h2f_loan_in[44] ),
	.h2f_loan_in_45(\hps_0|fpga_interfaces|h2f_loan_in[45] ),
	.h2f_loan_in_46(\hps_0|fpga_interfaces|h2f_loan_in[46] ),
	.h2f_loan_in_47(\hps_0|fpga_interfaces|h2f_loan_in[47] ),
	.h2f_loan_in_48(\hps_0|fpga_interfaces|h2f_loan_in[48] ),
	.h2f_loan_in_49(\hps_0|fpga_interfaces|h2f_loan_in[49] ),
	.h2f_loan_in_50(\hps_0|fpga_interfaces|h2f_loan_in[50] ),
	.h2f_loan_in_51(\hps_0|fpga_interfaces|h2f_loan_in[51] ),
	.h2f_loan_in_52(\hps_0|fpga_interfaces|h2f_loan_in[52] ),
	.h2f_loan_in_53(\hps_0|fpga_interfaces|h2f_loan_in[53] ),
	.h2f_loan_in_54(\hps_0|fpga_interfaces|h2f_loan_in[54] ),
	.h2f_loan_in_55(\hps_0|fpga_interfaces|h2f_loan_in[55] ),
	.h2f_loan_in_56(\hps_0|fpga_interfaces|h2f_loan_in[56] ),
	.h2f_loan_in_57(\hps_0|fpga_interfaces|h2f_loan_in[57] ),
	.h2f_loan_in_58(\hps_0|fpga_interfaces|h2f_loan_in[58] ),
	.h2f_loan_in_59(\hps_0|fpga_interfaces|h2f_loan_in[59] ),
	.h2f_loan_in_60(\hps_0|fpga_interfaces|h2f_loan_in[60] ),
	.h2f_loan_in_61(\hps_0|fpga_interfaces|h2f_loan_in[61] ),
	.h2f_loan_in_62(\hps_0|fpga_interfaces|h2f_loan_in[62] ),
	.h2f_loan_in_63(\hps_0|fpga_interfaces|h2f_loan_in[63] ),
	.h2f_loan_in_64(\hps_0|fpga_interfaces|h2f_loan_in[64] ),
	.h2f_loan_in_65(\hps_0|fpga_interfaces|h2f_loan_in[65] ),
	.h2f_loan_in_66(\hps_0|fpga_interfaces|h2f_loan_in[66] ),
	.h2f_rst_n_0(\hps_0|fpga_interfaces|h2f_rst_n[0] ),
	.h2f_lw_ARVALID_0(\hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps_0|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps_0|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps_0|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps_0|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\hps_0|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARADDR_6(\hps_0|fpga_interfaces|h2f_lw_ARADDR[6] ),
	.h2f_lw_ARADDR_7(\hps_0|fpga_interfaces|h2f_lw_ARADDR[7] ),
	.h2f_lw_ARADDR_8(\hps_0|fpga_interfaces|h2f_lw_ARADDR[8] ),
	.h2f_lw_ARADDR_9(\hps_0|fpga_interfaces|h2f_lw_ARADDR[9] ),
	.h2f_lw_ARADDR_10(\hps_0|fpga_interfaces|h2f_lw_ARADDR[10] ),
	.h2f_lw_ARADDR_11(\hps_0|fpga_interfaces|h2f_lw_ARADDR[11] ),
	.h2f_lw_ARADDR_12(\hps_0|fpga_interfaces|h2f_lw_ARADDR[12] ),
	.h2f_lw_ARADDR_13(\hps_0|fpga_interfaces|h2f_lw_ARADDR[13] ),
	.h2f_lw_ARADDR_14(\hps_0|fpga_interfaces|h2f_lw_ARADDR[14] ),
	.h2f_lw_ARBURST_0(\hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps_0|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps_0|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps_0|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps_0|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps_0|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps_0|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps_0|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps_0|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps_0|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps_0|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps_0|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps_0|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\hps_0|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWADDR_6(\hps_0|fpga_interfaces|h2f_lw_AWADDR[6] ),
	.h2f_lw_AWADDR_7(\hps_0|fpga_interfaces|h2f_lw_AWADDR[7] ),
	.h2f_lw_AWADDR_8(\hps_0|fpga_interfaces|h2f_lw_AWADDR[8] ),
	.h2f_lw_AWADDR_9(\hps_0|fpga_interfaces|h2f_lw_AWADDR[9] ),
	.h2f_lw_AWADDR_10(\hps_0|fpga_interfaces|h2f_lw_AWADDR[10] ),
	.h2f_lw_AWADDR_11(\hps_0|fpga_interfaces|h2f_lw_AWADDR[11] ),
	.h2f_lw_AWADDR_12(\hps_0|fpga_interfaces|h2f_lw_AWADDR[12] ),
	.h2f_lw_AWADDR_13(\hps_0|fpga_interfaces|h2f_lw_AWADDR[13] ),
	.h2f_lw_AWADDR_14(\hps_0|fpga_interfaces|h2f_lw_AWADDR[14] ),
	.h2f_lw_AWBURST_0(\hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps_0|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps_0|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps_0|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps_0|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps_0|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps_0|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps_0|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps_0|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps_0|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps_0|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps_0|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps_0|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps_0|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps_0|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps_0|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps_0|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps_0|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps_0|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps_0|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps_0|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps_0|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps_0|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps_0|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps_0|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps_0|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps_0|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps_0|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps_0|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps_0|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps_0|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps_0|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps_0|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps_0|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps_0|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps_0|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps_0|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps_0|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps_0|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps_0|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps_0|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps_0|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps_0|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps_0|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps_0|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.sink1_ready(\mm_interconnect_0|cmd_mux|sink1_ready~combout ),
	.awready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~combout ),
	.source_endofpacket(\mm_interconnect_0|onchip_memory2_0_s1_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.wready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_88_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][99]~q ),
	.out_data_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[7]~7_combout ),
	.out_data_8(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[8]~8_combout ),
	.out_data_9(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[9]~9_combout ),
	.out_data_10(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[10]~10_combout ),
	.out_data_11(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[11]~11_combout ),
	.out_data_12(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[12]~12_combout ),
	.out_data_13(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[13]~13_combout ),
	.out_data_14(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[14]~14_combout ),
	.out_data_15(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[15]~15_combout ),
	.out_data_16(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[16]~16_combout ),
	.out_data_17(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[17]~17_combout ),
	.out_data_18(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[18]~18_combout ),
	.out_data_19(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[19]~19_combout ),
	.out_data_20(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[20]~20_combout ),
	.out_data_21(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[21]~21_combout ),
	.out_data_22(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[22]~22_combout ),
	.out_data_23(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[23]~23_combout ),
	.out_data_24(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[24]~24_combout ),
	.out_data_25(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[25]~25_combout ),
	.out_data_26(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[26]~26_combout ),
	.out_data_27(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[27]~27_combout ),
	.out_data_28(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[28]~28_combout ),
	.out_data_29(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[29]~29_combout ),
	.out_data_30(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[30]~30_combout ),
	.out_data_31(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[31]~31_combout ),
	.emac1_inst(\hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ),
	.emac1_inst1(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ),
	.intermediate_0(\hps_0|hps_io|border|intermediate[0] ),
	.intermediate_1(\hps_0|hps_io|border|intermediate[1] ),
	.emac1_inst2(\hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ),
	.emac1_inst3(\hps_0|hps_io|border|emac1_inst~emac_phy_txd ),
	.emac1_inst4(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ),
	.emac1_inst5(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ),
	.emac1_inst6(\hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ),
	.qspi_inst(\hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ),
	.intermediate_2(\hps_0|hps_io|border|intermediate[2] ),
	.intermediate_4(\hps_0|hps_io|border|intermediate[4] ),
	.intermediate_6(\hps_0|hps_io|border|intermediate[6] ),
	.intermediate_8(\hps_0|hps_io|border|intermediate[8] ),
	.intermediate_3(\hps_0|hps_io|border|intermediate[3] ),
	.intermediate_5(\hps_0|hps_io|border|intermediate[5] ),
	.intermediate_7(\hps_0|hps_io|border|intermediate[7] ),
	.intermediate_9(\hps_0|hps_io|border|intermediate[9] ),
	.qspi_inst1(\hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ),
	.sdio_inst(\hps_0|hps_io|border|sdio_inst~sdmmc_cclk ),
	.intermediate_10(\hps_0|hps_io|border|intermediate[10] ),
	.intermediate_11(\hps_0|hps_io|border|intermediate[11] ),
	.intermediate_12(\hps_0|hps_io|border|intermediate[12] ),
	.intermediate_14(\hps_0|hps_io|border|intermediate[14] ),
	.intermediate_16(\hps_0|hps_io|border|intermediate[16] ),
	.intermediate_18(\hps_0|hps_io|border|intermediate[18] ),
	.intermediate_13(\hps_0|hps_io|border|intermediate[13] ),
	.intermediate_15(\hps_0|hps_io|border|intermediate[15] ),
	.intermediate_17(\hps_0|hps_io|border|intermediate[17] ),
	.intermediate_19(\hps_0|hps_io|border|intermediate[19] ),
	.usb1_inst(\hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ),
	.intermediate_20(\hps_0|hps_io|border|intermediate[20] ),
	.intermediate_22(\hps_0|hps_io|border|intermediate[22] ),
	.intermediate_24(\hps_0|hps_io|border|intermediate[24] ),
	.intermediate_26(\hps_0|hps_io|border|intermediate[26] ),
	.intermediate_28(\hps_0|hps_io|border|intermediate[28] ),
	.intermediate_30(\hps_0|hps_io|border|intermediate[30] ),
	.intermediate_32(\hps_0|hps_io|border|intermediate[32] ),
	.intermediate_34(\hps_0|hps_io|border|intermediate[34] ),
	.intermediate_21(\hps_0|hps_io|border|intermediate[21] ),
	.intermediate_23(\hps_0|hps_io|border|intermediate[23] ),
	.intermediate_25(\hps_0|hps_io|border|intermediate[25] ),
	.intermediate_27(\hps_0|hps_io|border|intermediate[27] ),
	.intermediate_29(\hps_0|hps_io|border|intermediate[29] ),
	.intermediate_31(\hps_0|hps_io|border|intermediate[31] ),
	.intermediate_33(\hps_0|hps_io|border|intermediate[33] ),
	.intermediate_35(\hps_0|hps_io|border|intermediate[35] ),
	.spim0_inst(\hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SCLK ),
	.spim0_inst1(\hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SS_0_N ),
	.intermediate_36(\hps_0|hps_io|border|intermediate[36] ),
	.intermediate_37(\hps_0|hps_io|border|intermediate[37] ),
	.spim1_inst(\hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ),
	.spim1_inst1(\hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ),
	.intermediate_38(\hps_0|hps_io|border|intermediate[38] ),
	.intermediate_39(\hps_0|hps_io|border|intermediate[39] ),
	.uart0_inst(\hps_0|hps_io|border|uart0_inst~uart_txd ),
	.intermediate_50(\hps_0|hps_io|border|intermediate[50] ),
	.intermediate_40(\hps_0|hps_io|border|intermediate[40] ),
	.intermediate_51(\hps_0|hps_io|border|intermediate[51] ),
	.intermediate_41(\hps_0|hps_io|border|intermediate[41] ),
	.intermediate_42(\hps_0|hps_io|border|intermediate[42] ),
	.intermediate_52(\hps_0|hps_io|border|intermediate[52] ),
	.intermediate_44(\hps_0|hps_io|border|intermediate[44] ),
	.intermediate_54(\hps_0|hps_io|border|intermediate[54] ),
	.intermediate_56(\hps_0|hps_io|border|intermediate[56] ),
	.intermediate_58(\hps_0|hps_io|border|intermediate[58] ),
	.intermediate_60(\hps_0|hps_io|border|intermediate[60] ),
	.intermediate_62(\hps_0|hps_io|border|intermediate[62] ),
	.intermediate_64(\hps_0|hps_io|border|intermediate[64] ),
	.intermediate_43(\hps_0|hps_io|border|intermediate[43] ),
	.intermediate_53(\hps_0|hps_io|border|intermediate[53] ),
	.intermediate_45(\hps_0|hps_io|border|intermediate[45] ),
	.intermediate_55(\hps_0|hps_io|border|intermediate[55] ),
	.intermediate_57(\hps_0|hps_io|border|intermediate[57] ),
	.intermediate_59(\hps_0|hps_io|border|intermediate[59] ),
	.intermediate_61(\hps_0|hps_io|border|intermediate[61] ),
	.intermediate_63(\hps_0|hps_io|border|intermediate[63] ),
	.intermediate_65(\hps_0|hps_io|border|intermediate[65] ),
	.intermediate_46(\hps_0|hps_io|border|intermediate[46] ),
	.intermediate_48(\hps_0|hps_io|border|intermediate[48] ),
	.intermediate_47(\hps_0|hps_io|border|intermediate[47] ),
	.intermediate_49(\hps_0|hps_io|border|intermediate[49] ),
	.parallelterminationcontrol_0(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ),
	.parallelterminationcontrol_1(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ),
	.parallelterminationcontrol_2(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ),
	.parallelterminationcontrol_3(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ),
	.parallelterminationcontrol_4(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ),
	.parallelterminationcontrol_5(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ),
	.parallelterminationcontrol_6(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ),
	.parallelterminationcontrol_7(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ),
	.parallelterminationcontrol_8(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ),
	.parallelterminationcontrol_9(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ),
	.parallelterminationcontrol_10(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ),
	.parallelterminationcontrol_11(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ),
	.parallelterminationcontrol_12(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ),
	.parallelterminationcontrol_13(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ),
	.parallelterminationcontrol_14(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ),
	.parallelterminationcontrol_15(\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ),
	.seriesterminationcontrol_0(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ),
	.seriesterminationcontrol_1(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ),
	.seriesterminationcontrol_2(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ),
	.seriesterminationcontrol_3(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ),
	.seriesterminationcontrol_4(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ),
	.seriesterminationcontrol_5(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ),
	.seriesterminationcontrol_6(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ),
	.seriesterminationcontrol_7(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ),
	.seriesterminationcontrol_8(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ),
	.seriesterminationcontrol_9(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ),
	.seriesterminationcontrol_10(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ),
	.seriesterminationcontrol_11(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ),
	.seriesterminationcontrol_12(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ),
	.seriesterminationcontrol_13(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ),
	.seriesterminationcontrol_14(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ),
	.seriesterminationcontrol_15(\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ),
	.dqsin(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dataout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ),
	.dataout_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ),
	.dataout_2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ),
	.dataout_3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ),
	.dataout_4(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ),
	.dataout_5(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ),
	.dataout_6(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ),
	.dataout_7(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ),
	.dataout_8(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ),
	.dataout_9(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ),
	.dataout_10(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ),
	.dataout_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ),
	.dataout_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ),
	.dataout_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ),
	.dataout_14(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ),
	.dataout_01(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ),
	.dataout_15(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ),
	.dataout_21(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ),
	.dataout_16(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ),
	.dataout_02(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ),
	.dataout_31(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ),
	.dataout_41(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ),
	.dataout_51(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ),
	.dataout_03(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ),
	.dataout_22(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ),
	.extra_output_pad_gen0delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.wire_pseudo_diffa_o_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.wire_pseudo_diffa_obar_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.wire_pseudo_diffa_oeout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.wire_pseudo_diffa_oebout_0(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.pad_gen0delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_11(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_12(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_13(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.os(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar1(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar2(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar3(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.hps_io_emac1_inst_MDIO_0(\hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ),
	.hps_io_qspi_inst_IO0_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ),
	.hps_io_qspi_inst_IO1_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ),
	.hps_io_qspi_inst_IO2_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ),
	.hps_io_qspi_inst_IO3_0(\hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ),
	.hps_io_sdio_inst_CMD_0(\hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ),
	.hps_io_sdio_inst_D0_0(\hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ),
	.hps_io_sdio_inst_D1_0(\hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ),
	.hps_io_sdio_inst_D2_0(\hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ),
	.hps_io_sdio_inst_D3_0(\hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D0_0(\hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ),
	.hps_io_usb1_inst_D1_0(\hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ),
	.hps_io_usb1_inst_D2_0(\hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ),
	.hps_io_usb1_inst_D3_0(\hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D4_0(\hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ),
	.hps_io_usb1_inst_D5_0(\hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ),
	.hps_io_usb1_inst_D6_0(\hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ),
	.hps_io_usb1_inst_D7_0(\hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ),
	.hps_io_gpio_inst_GPIO09_0(\hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ),
	.hps_io_gpio_inst_GPIO40_0(\hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ),
	.hps_io_gpio_inst_GPIO48_0(\hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ),
	.hps_io_gpio_inst_GPIO61_0(\hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ),
	.hps_io_gpio_inst_GPIO62_0(\hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~input_o ),
	.hps_io_gpio_inst_LOANIO00_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~input_o ),
	.hps_io_gpio_inst_LOANIO41_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~input_o ),
	.hps_io_gpio_inst_LOANIO51_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~input_o ),
	.hps_io_gpio_inst_LOANIO52_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~input_o ),
	.hps_io_gpio_inst_LOANIO53_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~input_o ),
	.hps_io_gpio_inst_LOANIO54_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~input_o ),
	.hps_io_gpio_inst_LOANIO55_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~input_o ),
	.hps_io_gpio_inst_LOANIO56_0(\hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~input_o ),
	.hps_io_hps_io_emac1_inst_RXD0(\hps_io_hps_io_emac1_inst_RXD0~input_o ),
	.hps_io_hps_io_emac1_inst_RXD1(\hps_io_hps_io_emac1_inst_RXD1~input_o ),
	.hps_io_hps_io_emac1_inst_RXD2(\hps_io_hps_io_emac1_inst_RXD2~input_o ),
	.hps_io_hps_io_emac1_inst_RXD3(\hps_io_hps_io_emac1_inst_RXD3~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CLK(\hps_io_hps_io_emac1_inst_RX_CLK~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CTL(\hps_io_hps_io_emac1_inst_RX_CTL~input_o ),
	.hps_io_hps_io_spim0_inst_MISO(\hps_io_hps_io_spim0_inst_MISO~input_o ),
	.hps_io_hps_io_spim1_inst_MISO(\hps_io_hps_io_spim1_inst_MISO~input_o ),
	.hps_io_hps_io_uart0_inst_RX(\hps_io_hps_io_uart0_inst_RX~input_o ),
	.hps_io_hps_io_usb1_inst_CLK(\hps_io_hps_io_usb1_inst_CLK~input_o ),
	.hps_io_hps_io_usb1_inst_DIR(\hps_io_hps_io_usb1_inst_DIR~input_o ),
	.hps_io_hps_io_usb1_inst_NXT(\hps_io_hps_io_usb1_inst_NXT~input_o ),
	.memory_oct_rzqin(\memory_oct_rzqin~input_o ),
	.d_out_oe_0(\d_out_oe[0]~input_o ),
	.d_out_oe_1(\d_out_oe[1]~input_o ),
	.d_out_oe_2(\d_out_oe[2]~input_o ),
	.d_out_oe_3(\d_out_oe[3]~input_o ),
	.d_out_oe_4(\d_out_oe[4]~input_o ),
	.d_out_oe_5(\d_out_oe[5]~input_o ),
	.d_out_oe_6(\d_out_oe[6]~input_o ),
	.d_out_oe_7(\d_out_oe[7]~input_o ),
	.d_out_oe_8(\d_out_oe[8]~input_o ),
	.d_out_oe_9(\d_out_oe[9]~input_o ),
	.d_out_oe_10(\d_out_oe[10]~input_o ),
	.d_out_oe_11(\d_out_oe[11]~input_o ),
	.d_out_oe_12(\d_out_oe[12]~input_o ),
	.d_out_oe_13(\d_out_oe[13]~input_o ),
	.d_out_oe_14(\d_out_oe[14]~input_o ),
	.d_out_oe_15(\d_out_oe[15]~input_o ),
	.d_out_oe_16(\d_out_oe[16]~input_o ),
	.d_out_oe_17(\d_out_oe[17]~input_o ),
	.d_out_oe_18(\d_out_oe[18]~input_o ),
	.d_out_oe_19(\d_out_oe[19]~input_o ),
	.d_out_oe_20(\d_out_oe[20]~input_o ),
	.d_out_oe_21(\d_out_oe[21]~input_o ),
	.d_out_oe_22(\d_out_oe[22]~input_o ),
	.d_out_oe_23(\d_out_oe[23]~input_o ),
	.d_out_oe_24(\d_out_oe[24]~input_o ),
	.d_out_oe_25(\d_out_oe[25]~input_o ),
	.d_out_oe_26(\d_out_oe[26]~input_o ),
	.d_out_oe_27(\d_out_oe[27]~input_o ),
	.d_out_oe_28(\d_out_oe[28]~input_o ),
	.d_out_oe_29(\d_out_oe[29]~input_o ),
	.d_out_oe_30(\d_out_oe[30]~input_o ),
	.d_out_oe_31(\d_out_oe[31]~input_o ),
	.d_out_oe_32(\d_out_oe[32]~input_o ),
	.d_out_oe_33(\d_out_oe[33]~input_o ),
	.d_out_oe_34(\d_out_oe[34]~input_o ),
	.d_out_oe_35(\d_out_oe[35]~input_o ),
	.d_out_oe_36(\d_out_oe[36]~input_o ),
	.d_out_oe_37(\d_out_oe[37]~input_o ),
	.d_out_oe_38(\d_out_oe[38]~input_o ),
	.d_out_oe_39(\d_out_oe[39]~input_o ),
	.d_out_oe_40(\d_out_oe[40]~input_o ),
	.d_out_oe_41(\d_out_oe[41]~input_o ),
	.d_out_oe_42(\d_out_oe[42]~input_o ),
	.d_out_oe_43(\d_out_oe[43]~input_o ),
	.d_out_oe_44(\d_out_oe[44]~input_o ),
	.d_out_oe_45(\d_out_oe[45]~input_o ),
	.d_out_oe_46(\d_out_oe[46]~input_o ),
	.d_out_oe_47(\d_out_oe[47]~input_o ),
	.d_out_oe_48(\d_out_oe[48]~input_o ),
	.d_out_oe_49(\d_out_oe[49]~input_o ),
	.d_out_oe_50(\d_out_oe[50]~input_o ),
	.d_out_oe_51(\d_out_oe[51]~input_o ),
	.d_out_oe_52(\d_out_oe[52]~input_o ),
	.d_out_oe_53(\d_out_oe[53]~input_o ),
	.d_out_oe_54(\d_out_oe[54]~input_o ),
	.d_out_oe_55(\d_out_oe[55]~input_o ),
	.d_out_oe_56(\d_out_oe[56]~input_o ),
	.d_out_oe_57(\d_out_oe[57]~input_o ),
	.d_out_oe_58(\d_out_oe[58]~input_o ),
	.d_out_oe_59(\d_out_oe[59]~input_o ),
	.d_out_oe_60(\d_out_oe[60]~input_o ),
	.d_out_oe_61(\d_out_oe[61]~input_o ),
	.d_out_oe_62(\d_out_oe[62]~input_o ),
	.d_out_oe_63(\d_out_oe[63]~input_o ),
	.d_out_oe_64(\d_out_oe[64]~input_o ),
	.d_out_oe_65(\d_out_oe[65]~input_o ),
	.d_out_oe_66(\d_out_oe[66]~input_o ),
	.d_out_out_0(\d_out_out[0]~input_o ),
	.d_out_out_1(\d_out_out[1]~input_o ),
	.d_out_out_2(\d_out_out[2]~input_o ),
	.d_out_out_3(\d_out_out[3]~input_o ),
	.d_out_out_4(\d_out_out[4]~input_o ),
	.d_out_out_5(\d_out_out[5]~input_o ),
	.d_out_out_6(\d_out_out[6]~input_o ),
	.d_out_out_7(\d_out_out[7]~input_o ),
	.d_out_out_8(\d_out_out[8]~input_o ),
	.d_out_out_9(\d_out_out[9]~input_o ),
	.d_out_out_10(\d_out_out[10]~input_o ),
	.d_out_out_11(\d_out_out[11]~input_o ),
	.d_out_out_12(\d_out_out[12]~input_o ),
	.d_out_out_13(\d_out_out[13]~input_o ),
	.d_out_out_14(\d_out_out[14]~input_o ),
	.d_out_out_15(\d_out_out[15]~input_o ),
	.d_out_out_16(\d_out_out[16]~input_o ),
	.d_out_out_17(\d_out_out[17]~input_o ),
	.d_out_out_18(\d_out_out[18]~input_o ),
	.d_out_out_19(\d_out_out[19]~input_o ),
	.d_out_out_20(\d_out_out[20]~input_o ),
	.d_out_out_21(\d_out_out[21]~input_o ),
	.d_out_out_22(\d_out_out[22]~input_o ),
	.d_out_out_23(\d_out_out[23]~input_o ),
	.d_out_out_24(\d_out_out[24]~input_o ),
	.d_out_out_25(\d_out_out[25]~input_o ),
	.d_out_out_26(\d_out_out[26]~input_o ),
	.d_out_out_27(\d_out_out[27]~input_o ),
	.d_out_out_28(\d_out_out[28]~input_o ),
	.d_out_out_29(\d_out_out[29]~input_o ),
	.d_out_out_30(\d_out_out[30]~input_o ),
	.d_out_out_31(\d_out_out[31]~input_o ),
	.d_out_out_32(\d_out_out[32]~input_o ),
	.d_out_out_33(\d_out_out[33]~input_o ),
	.d_out_out_34(\d_out_out[34]~input_o ),
	.d_out_out_35(\d_out_out[35]~input_o ),
	.d_out_out_36(\d_out_out[36]~input_o ),
	.d_out_out_37(\d_out_out[37]~input_o ),
	.d_out_out_38(\d_out_out[38]~input_o ),
	.d_out_out_39(\d_out_out[39]~input_o ),
	.d_out_out_40(\d_out_out[40]~input_o ),
	.d_out_out_41(\d_out_out[41]~input_o ),
	.d_out_out_42(\d_out_out[42]~input_o ),
	.d_out_out_43(\d_out_out[43]~input_o ),
	.d_out_out_44(\d_out_out[44]~input_o ),
	.d_out_out_45(\d_out_out[45]~input_o ),
	.d_out_out_46(\d_out_out[46]~input_o ),
	.d_out_out_47(\d_out_out[47]~input_o ),
	.d_out_out_48(\d_out_out[48]~input_o ),
	.d_out_out_49(\d_out_out[49]~input_o ),
	.d_out_out_50(\d_out_out[50]~input_o ),
	.d_out_out_51(\d_out_out[51]~input_o ),
	.d_out_out_52(\d_out_out[52]~input_o ),
	.d_out_out_53(\d_out_out[53]~input_o ),
	.d_out_out_54(\d_out_out[54]~input_o ),
	.d_out_out_55(\d_out_out[55]~input_o ),
	.d_out_out_56(\d_out_out[56]~input_o ),
	.d_out_out_57(\d_out_out[57]~input_o ),
	.d_out_out_58(\d_out_out[58]~input_o ),
	.d_out_out_59(\d_out_out[59]~input_o ),
	.d_out_out_60(\d_out_out[60]~input_o ),
	.d_out_out_61(\d_out_out[61]~input_o ),
	.d_out_out_62(\d_out_out[62]~input_o ),
	.d_out_out_63(\d_out_out[63]~input_o ),
	.d_out_out_64(\d_out_out[64]~input_o ),
	.d_out_out_65(\d_out_out[65]~input_o ),
	.d_out_out_66(\d_out_out[66]~input_o ));

soc_system_soc_system_mm_interconnect_0 mm_interconnect_0(
	.h2f_lw_ARVALID_0(\hps_0|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps_0|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps_0|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps_0|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps_0|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps_0|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps_0|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps_0|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps_0|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps_0|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps_0|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\hps_0|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARADDR_6(\hps_0|fpga_interfaces|h2f_lw_ARADDR[6] ),
	.h2f_lw_ARADDR_7(\hps_0|fpga_interfaces|h2f_lw_ARADDR[7] ),
	.h2f_lw_ARADDR_8(\hps_0|fpga_interfaces|h2f_lw_ARADDR[8] ),
	.h2f_lw_ARADDR_9(\hps_0|fpga_interfaces|h2f_lw_ARADDR[9] ),
	.h2f_lw_ARADDR_10(\hps_0|fpga_interfaces|h2f_lw_ARADDR[10] ),
	.h2f_lw_ARADDR_11(\hps_0|fpga_interfaces|h2f_lw_ARADDR[11] ),
	.h2f_lw_ARADDR_12(\hps_0|fpga_interfaces|h2f_lw_ARADDR[12] ),
	.h2f_lw_ARADDR_13(\hps_0|fpga_interfaces|h2f_lw_ARADDR[13] ),
	.h2f_lw_ARADDR_14(\hps_0|fpga_interfaces|h2f_lw_ARADDR[14] ),
	.h2f_lw_ARBURST_0(\hps_0|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps_0|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps_0|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps_0|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps_0|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps_0|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps_0|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps_0|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps_0|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps_0|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps_0|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps_0|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps_0|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps_0|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps_0|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps_0|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps_0|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps_0|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps_0|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps_0|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps_0|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps_0|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps_0|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps_0|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\hps_0|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWADDR_6(\hps_0|fpga_interfaces|h2f_lw_AWADDR[6] ),
	.h2f_lw_AWADDR_7(\hps_0|fpga_interfaces|h2f_lw_AWADDR[7] ),
	.h2f_lw_AWADDR_8(\hps_0|fpga_interfaces|h2f_lw_AWADDR[8] ),
	.h2f_lw_AWADDR_9(\hps_0|fpga_interfaces|h2f_lw_AWADDR[9] ),
	.h2f_lw_AWADDR_10(\hps_0|fpga_interfaces|h2f_lw_AWADDR[10] ),
	.h2f_lw_AWADDR_11(\hps_0|fpga_interfaces|h2f_lw_AWADDR[11] ),
	.h2f_lw_AWADDR_12(\hps_0|fpga_interfaces|h2f_lw_AWADDR[12] ),
	.h2f_lw_AWADDR_13(\hps_0|fpga_interfaces|h2f_lw_AWADDR[13] ),
	.h2f_lw_AWADDR_14(\hps_0|fpga_interfaces|h2f_lw_AWADDR[14] ),
	.h2f_lw_AWBURST_0(\hps_0|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps_0|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps_0|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps_0|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps_0|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps_0|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps_0|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps_0|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps_0|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps_0|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps_0|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps_0|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps_0|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps_0|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps_0|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps_0|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps_0|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps_0|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps_0|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps_0|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps_0|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps_0|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps_0|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps_0|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps_0|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps_0|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps_0|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps_0|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps_0|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps_0|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps_0|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps_0|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps_0|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps_0|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps_0|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps_0|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps_0|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps_0|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps_0|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps_0|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps_0|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps_0|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps_0|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps_0|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps_0|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps_0|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps_0|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps_0|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps_0|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps_0|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps_0|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps_0|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps_0|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps_0|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps_0|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.source0_data_34(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~2_combout ),
	.source0_data_32(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~3_combout ),
	.sink1_ready(\mm_interconnect_0|cmd_mux|sink1_ready~combout ),
	.hps_0_h2f_lw_axi_master_awready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux|src0_valid~combout ),
	.source_endofpacket(\mm_interconnect_0|onchip_memory2_0_s1_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_0|rsp_demux|src1_valid~0_combout ),
	.hps_0_h2f_lw_axi_master_wready(\mm_interconnect_0|hps_0_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_88_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem[0][99]~q ),
	.out_data_0(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[7]~7_combout ),
	.out_data_8(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[8]~8_combout ),
	.out_data_9(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[9]~9_combout ),
	.out_data_10(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[10]~10_combout ),
	.out_data_11(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[11]~11_combout ),
	.out_data_12(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[12]~12_combout ),
	.out_data_13(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[13]~13_combout ),
	.out_data_14(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[14]~14_combout ),
	.out_data_15(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[15]~15_combout ),
	.out_data_16(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[16]~16_combout ),
	.out_data_17(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[17]~17_combout ),
	.out_data_18(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[18]~18_combout ),
	.out_data_19(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[19]~19_combout ),
	.out_data_20(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[20]~20_combout ),
	.out_data_21(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[21]~21_combout ),
	.out_data_22(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[22]~22_combout ),
	.out_data_23(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[23]~23_combout ),
	.out_data_24(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[24]~24_combout ),
	.out_data_25(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[25]~25_combout ),
	.out_data_26(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[26]~26_combout ),
	.out_data_27(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[27]~27_combout ),
	.out_data_28(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[28]~28_combout ),
	.out_data_29(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[29]~29_combout ),
	.out_data_30(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[30]~30_combout ),
	.out_data_31(\mm_interconnect_0|onchip_memory2_0_s1_agent_rdata_fifo|out_data[31]~31_combout ),
	.m0_write(\mm_interconnect_0|onchip_memory2_0_s1_agent|m0_write~1_combout ),
	.in_data_reg_0(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_5(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ),
	.int_nxt_addr_reg_dly_6(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ),
	.int_nxt_addr_reg_dly_7(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ),
	.int_nxt_addr_reg_dly_8(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ),
	.int_nxt_addr_reg_dly_9(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ),
	.int_nxt_addr_reg_dly_10(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[10]~q ),
	.int_nxt_addr_reg_dly_11(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[11]~q ),
	.int_nxt_addr_reg_dly_12(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[12]~q ),
	.int_nxt_addr_reg_dly_13(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[13]~q ),
	.int_nxt_addr_reg_dly_14(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[14]~q ),
	.in_data_reg_1(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.source0_data_33(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~7_combout ),
	.in_data_reg_9(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.source0_data_35(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~8_combout ),
	.in_data_reg_25(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out1(\rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

soc_system_soc_system_pll_0 pll_0(
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

soc_system_soc_system_onchip_memory2_0 onchip_memory2_0(
	.outclk_wire_0(\pll_0|altera_pll_i|outclk_wire[0] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_b_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[0] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_b_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[1] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_b_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_b_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_b_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[4] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_b_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[5] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_b_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[6] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_b_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[7] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_b_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[8] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_b_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[9] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_b_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[10] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_b_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[11] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_b_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[12] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_b_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[13] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_b_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_b_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[15] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_b_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[16] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_b_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[17] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_b_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[18] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_b_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[19] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_b_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[20] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_b_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[21] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_b_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_b_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_b_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_b_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_b_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[26] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_b_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_b_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_b_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_b_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_b_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_b[31] ),
	.source0_data_34(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~2_combout ),
	.source0_data_32(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~3_combout ),
	.m0_write(\mm_interconnect_0|onchip_memory2_0_s1_agent|m0_write~1_combout ),
	.in_data_reg_0(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_5(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ),
	.int_nxt_addr_reg_dly_6(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ),
	.int_nxt_addr_reg_dly_7(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ),
	.int_nxt_addr_reg_dly_8(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ),
	.int_nxt_addr_reg_dly_9(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ),
	.int_nxt_addr_reg_dly_10(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[10]~q ),
	.int_nxt_addr_reg_dly_11(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[11]~q ),
	.int_nxt_addr_reg_dly_12(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[12]~q ),
	.int_nxt_addr_reg_dly_13(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[13]~q ),
	.int_nxt_addr_reg_dly_14(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[14]~q ),
	.in_data_reg_1(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.source0_data_33(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~7_combout ),
	.in_data_reg_9(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.source0_data_35(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~8_combout ),
	.in_data_reg_25(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.ram_mm_chipselect(\ram_mm_chipselect~input_o ),
	.ram_mm_write(\ram_mm_write~input_o ),
	.ram_clk_clk(\ram_clk_clk~input_o ),
	.ram_mm_clken(\ram_mm_clken~input_o ),
	.ram_mm_writedata_0(\ram_mm_writedata[0]~input_o ),
	.ram_mm_address_0(\ram_mm_address[0]~input_o ),
	.ram_mm_address_1(\ram_mm_address[1]~input_o ),
	.ram_mm_address_2(\ram_mm_address[2]~input_o ),
	.ram_mm_address_3(\ram_mm_address[3]~input_o ),
	.ram_mm_address_4(\ram_mm_address[4]~input_o ),
	.ram_mm_address_5(\ram_mm_address[5]~input_o ),
	.ram_mm_address_6(\ram_mm_address[6]~input_o ),
	.ram_mm_address_7(\ram_mm_address[7]~input_o ),
	.ram_mm_address_8(\ram_mm_address[8]~input_o ),
	.ram_mm_address_9(\ram_mm_address[9]~input_o ),
	.ram_mm_address_10(\ram_mm_address[10]~input_o ),
	.ram_mm_address_11(\ram_mm_address[11]~input_o ),
	.ram_mm_address_12(\ram_mm_address[12]~input_o ),
	.ram_mm_byteenable_0(\ram_mm_byteenable[0]~input_o ),
	.ram_mm_writedata_1(\ram_mm_writedata[1]~input_o ),
	.ram_mm_writedata_2(\ram_mm_writedata[2]~input_o ),
	.ram_mm_writedata_3(\ram_mm_writedata[3]~input_o ),
	.ram_mm_writedata_4(\ram_mm_writedata[4]~input_o ),
	.ram_mm_writedata_5(\ram_mm_writedata[5]~input_o ),
	.ram_mm_writedata_6(\ram_mm_writedata[6]~input_o ),
	.ram_mm_writedata_7(\ram_mm_writedata[7]~input_o ),
	.ram_mm_writedata_8(\ram_mm_writedata[8]~input_o ),
	.ram_mm_byteenable_1(\ram_mm_byteenable[1]~input_o ),
	.ram_mm_writedata_9(\ram_mm_writedata[9]~input_o ),
	.ram_mm_writedata_10(\ram_mm_writedata[10]~input_o ),
	.ram_mm_writedata_11(\ram_mm_writedata[11]~input_o ),
	.ram_mm_writedata_12(\ram_mm_writedata[12]~input_o ),
	.ram_mm_writedata_13(\ram_mm_writedata[13]~input_o ),
	.ram_mm_writedata_14(\ram_mm_writedata[14]~input_o ),
	.ram_mm_writedata_15(\ram_mm_writedata[15]~input_o ),
	.ram_mm_writedata_16(\ram_mm_writedata[16]~input_o ),
	.ram_mm_byteenable_2(\ram_mm_byteenable[2]~input_o ),
	.ram_mm_writedata_17(\ram_mm_writedata[17]~input_o ),
	.ram_mm_writedata_18(\ram_mm_writedata[18]~input_o ),
	.ram_mm_writedata_19(\ram_mm_writedata[19]~input_o ),
	.ram_mm_writedata_20(\ram_mm_writedata[20]~input_o ),
	.ram_mm_writedata_21(\ram_mm_writedata[21]~input_o ),
	.ram_mm_writedata_22(\ram_mm_writedata[22]~input_o ),
	.ram_mm_writedata_23(\ram_mm_writedata[23]~input_o ),
	.ram_mm_writedata_24(\ram_mm_writedata[24]~input_o ),
	.ram_mm_byteenable_3(\ram_mm_byteenable[3]~input_o ),
	.ram_mm_writedata_25(\ram_mm_writedata[25]~input_o ),
	.ram_mm_writedata_26(\ram_mm_writedata[26]~input_o ),
	.ram_mm_writedata_27(\ram_mm_writedata[27]~input_o ),
	.ram_mm_writedata_28(\ram_mm_writedata[28]~input_o ),
	.ram_mm_writedata_29(\ram_mm_writedata[29]~input_o ),
	.ram_mm_writedata_30(\ram_mm_writedata[30]~input_o ),
	.ram_mm_writedata_31(\ram_mm_writedata[31]~input_o ));

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[3]),
	.ibar(memory_mem_dqs_n[3]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[24]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[25]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[26]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[27]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[28]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[29]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[30]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[31]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[2]),
	.ibar(memory_mem_dqs_n[2]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[16]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[17]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[18]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[19]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[20]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[21]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[22]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[23]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[1]),
	.ibar(memory_mem_dqs_n[1]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[8]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[9]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[10]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[11]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[12]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[13]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[14]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[15]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[0]),
	.ibar(memory_mem_dqs_n[0]),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[0]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[1]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[2]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[3]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[4]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[5]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[6]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[7]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

assign \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o  = hps_io_hps_io_emac1_inst_MDIO;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o  = hps_io_hps_io_qspi_inst_IO0;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o  = hps_io_hps_io_qspi_inst_IO1;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o  = hps_io_hps_io_qspi_inst_IO2;

assign \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o  = hps_io_hps_io_qspi_inst_IO3;

assign \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o  = hps_io_hps_io_sdio_inst_CMD;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~input_o  = hps_io_hps_io_sdio_inst_D0;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~input_o  = hps_io_hps_io_sdio_inst_D1;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~input_o  = hps_io_hps_io_sdio_inst_D2;

assign \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~input_o  = hps_io_hps_io_sdio_inst_D3;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~input_o  = hps_io_hps_io_usb1_inst_D0;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~input_o  = hps_io_hps_io_usb1_inst_D1;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~input_o  = hps_io_hps_io_usb1_inst_D2;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~input_o  = hps_io_hps_io_usb1_inst_D3;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~input_o  = hps_io_hps_io_usb1_inst_D4;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~input_o  = hps_io_hps_io_usb1_inst_D5;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~input_o  = hps_io_hps_io_usb1_inst_D6;

assign \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~input_o  = hps_io_hps_io_usb1_inst_D7;

assign \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO09;

assign \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO40;

assign \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO48;

assign \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO61;

assign \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO62;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO00;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO41;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO51;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO52;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO53;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO54;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO55;

assign \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~input_o  = hps_io_hps_io_gpio_inst_LOANIO56;

assign \hps_io_hps_io_emac1_inst_RXD0~input_o  = hps_io_hps_io_emac1_inst_RXD0;

assign \hps_io_hps_io_emac1_inst_RXD1~input_o  = hps_io_hps_io_emac1_inst_RXD1;

assign \hps_io_hps_io_emac1_inst_RXD2~input_o  = hps_io_hps_io_emac1_inst_RXD2;

assign \hps_io_hps_io_emac1_inst_RXD3~input_o  = hps_io_hps_io_emac1_inst_RXD3;

assign \hps_io_hps_io_emac1_inst_RX_CLK~input_o  = hps_io_hps_io_emac1_inst_RX_CLK;

assign \hps_io_hps_io_emac1_inst_RX_CTL~input_o  = hps_io_hps_io_emac1_inst_RX_CTL;

assign \hps_io_hps_io_spim0_inst_MISO~input_o  = hps_io_hps_io_spim0_inst_MISO;

assign \hps_io_hps_io_spim1_inst_MISO~input_o  = hps_io_hps_io_spim1_inst_MISO;

assign \hps_io_hps_io_uart0_inst_RX~input_o  = hps_io_hps_io_uart0_inst_RX;

assign \hps_io_hps_io_usb1_inst_CLK~input_o  = hps_io_hps_io_usb1_inst_CLK;

assign \hps_io_hps_io_usb1_inst_DIR~input_o  = hps_io_hps_io_usb1_inst_DIR;

assign \hps_io_hps_io_usb1_inst_NXT~input_o  = hps_io_hps_io_usb1_inst_NXT;

assign \memory_oct_rzqin~input_o  = memory_oct_rzqin;

assign \d_out_oe[0]~input_o  = d_out_oe[0];

assign \d_out_oe[1]~input_o  = d_out_oe[1];

assign \d_out_oe[2]~input_o  = d_out_oe[2];

assign \d_out_oe[3]~input_o  = d_out_oe[3];

assign \d_out_oe[4]~input_o  = d_out_oe[4];

assign \d_out_oe[5]~input_o  = d_out_oe[5];

assign \d_out_oe[6]~input_o  = d_out_oe[6];

assign \d_out_oe[7]~input_o  = d_out_oe[7];

assign \d_out_oe[8]~input_o  = d_out_oe[8];

assign \d_out_oe[9]~input_o  = d_out_oe[9];

assign \d_out_oe[10]~input_o  = d_out_oe[10];

assign \d_out_oe[11]~input_o  = d_out_oe[11];

assign \d_out_oe[12]~input_o  = d_out_oe[12];

assign \d_out_oe[13]~input_o  = d_out_oe[13];

assign \d_out_oe[14]~input_o  = d_out_oe[14];

assign \d_out_oe[15]~input_o  = d_out_oe[15];

assign \d_out_oe[16]~input_o  = d_out_oe[16];

assign \d_out_oe[17]~input_o  = d_out_oe[17];

assign \d_out_oe[18]~input_o  = d_out_oe[18];

assign \d_out_oe[19]~input_o  = d_out_oe[19];

assign \d_out_oe[20]~input_o  = d_out_oe[20];

assign \d_out_oe[21]~input_o  = d_out_oe[21];

assign \d_out_oe[22]~input_o  = d_out_oe[22];

assign \d_out_oe[23]~input_o  = d_out_oe[23];

assign \d_out_oe[24]~input_o  = d_out_oe[24];

assign \d_out_oe[25]~input_o  = d_out_oe[25];

assign \d_out_oe[26]~input_o  = d_out_oe[26];

assign \d_out_oe[27]~input_o  = d_out_oe[27];

assign \d_out_oe[28]~input_o  = d_out_oe[28];

assign \d_out_oe[29]~input_o  = d_out_oe[29];

assign \d_out_oe[30]~input_o  = d_out_oe[30];

assign \d_out_oe[31]~input_o  = d_out_oe[31];

assign \d_out_oe[32]~input_o  = d_out_oe[32];

assign \d_out_oe[33]~input_o  = d_out_oe[33];

assign \d_out_oe[34]~input_o  = d_out_oe[34];

assign \d_out_oe[35]~input_o  = d_out_oe[35];

assign \d_out_oe[36]~input_o  = d_out_oe[36];

assign \d_out_oe[37]~input_o  = d_out_oe[37];

assign \d_out_oe[38]~input_o  = d_out_oe[38];

assign \d_out_oe[39]~input_o  = d_out_oe[39];

assign \d_out_oe[40]~input_o  = d_out_oe[40];

assign \d_out_oe[41]~input_o  = d_out_oe[41];

assign \d_out_oe[42]~input_o  = d_out_oe[42];

assign \d_out_oe[43]~input_o  = d_out_oe[43];

assign \d_out_oe[44]~input_o  = d_out_oe[44];

assign \d_out_oe[45]~input_o  = d_out_oe[45];

assign \d_out_oe[46]~input_o  = d_out_oe[46];

assign \d_out_oe[47]~input_o  = d_out_oe[47];

assign \d_out_oe[48]~input_o  = d_out_oe[48];

assign \d_out_oe[49]~input_o  = d_out_oe[49];

assign \d_out_oe[50]~input_o  = d_out_oe[50];

assign \d_out_oe[51]~input_o  = d_out_oe[51];

assign \d_out_oe[52]~input_o  = d_out_oe[52];

assign \d_out_oe[53]~input_o  = d_out_oe[53];

assign \d_out_oe[54]~input_o  = d_out_oe[54];

assign \d_out_oe[55]~input_o  = d_out_oe[55];

assign \d_out_oe[56]~input_o  = d_out_oe[56];

assign \d_out_oe[57]~input_o  = d_out_oe[57];

assign \d_out_oe[58]~input_o  = d_out_oe[58];

assign \d_out_oe[59]~input_o  = d_out_oe[59];

assign \d_out_oe[60]~input_o  = d_out_oe[60];

assign \d_out_oe[61]~input_o  = d_out_oe[61];

assign \d_out_oe[62]~input_o  = d_out_oe[62];

assign \d_out_oe[63]~input_o  = d_out_oe[63];

assign \d_out_oe[64]~input_o  = d_out_oe[64];

assign \d_out_oe[65]~input_o  = d_out_oe[65];

assign \d_out_oe[66]~input_o  = d_out_oe[66];

assign \d_out_out[0]~input_o  = d_out_out[0];

assign \d_out_out[1]~input_o  = d_out_out[1];

assign \d_out_out[2]~input_o  = d_out_out[2];

assign \d_out_out[3]~input_o  = d_out_out[3];

assign \d_out_out[4]~input_o  = d_out_out[4];

assign \d_out_out[5]~input_o  = d_out_out[5];

assign \d_out_out[6]~input_o  = d_out_out[6];

assign \d_out_out[7]~input_o  = d_out_out[7];

assign \d_out_out[8]~input_o  = d_out_out[8];

assign \d_out_out[9]~input_o  = d_out_out[9];

assign \d_out_out[10]~input_o  = d_out_out[10];

assign \d_out_out[11]~input_o  = d_out_out[11];

assign \d_out_out[12]~input_o  = d_out_out[12];

assign \d_out_out[13]~input_o  = d_out_out[13];

assign \d_out_out[14]~input_o  = d_out_out[14];

assign \d_out_out[15]~input_o  = d_out_out[15];

assign \d_out_out[16]~input_o  = d_out_out[16];

assign \d_out_out[17]~input_o  = d_out_out[17];

assign \d_out_out[18]~input_o  = d_out_out[18];

assign \d_out_out[19]~input_o  = d_out_out[19];

assign \d_out_out[20]~input_o  = d_out_out[20];

assign \d_out_out[21]~input_o  = d_out_out[21];

assign \d_out_out[22]~input_o  = d_out_out[22];

assign \d_out_out[23]~input_o  = d_out_out[23];

assign \d_out_out[24]~input_o  = d_out_out[24];

assign \d_out_out[25]~input_o  = d_out_out[25];

assign \d_out_out[26]~input_o  = d_out_out[26];

assign \d_out_out[27]~input_o  = d_out_out[27];

assign \d_out_out[28]~input_o  = d_out_out[28];

assign \d_out_out[29]~input_o  = d_out_out[29];

assign \d_out_out[30]~input_o  = d_out_out[30];

assign \d_out_out[31]~input_o  = d_out_out[31];

assign \d_out_out[32]~input_o  = d_out_out[32];

assign \d_out_out[33]~input_o  = d_out_out[33];

assign \d_out_out[34]~input_o  = d_out_out[34];

assign \d_out_out[35]~input_o  = d_out_out[35];

assign \d_out_out[36]~input_o  = d_out_out[36];

assign \d_out_out[37]~input_o  = d_out_out[37];

assign \d_out_out[38]~input_o  = d_out_out[38];

assign \d_out_out[39]~input_o  = d_out_out[39];

assign \d_out_out[40]~input_o  = d_out_out[40];

assign \d_out_out[41]~input_o  = d_out_out[41];

assign \d_out_out[42]~input_o  = d_out_out[42];

assign \d_out_out[43]~input_o  = d_out_out[43];

assign \d_out_out[44]~input_o  = d_out_out[44];

assign \d_out_out[45]~input_o  = d_out_out[45];

assign \d_out_out[46]~input_o  = d_out_out[46];

assign \d_out_out[47]~input_o  = d_out_out[47];

assign \d_out_out[48]~input_o  = d_out_out[48];

assign \d_out_out[49]~input_o  = d_out_out[49];

assign \d_out_out[50]~input_o  = d_out_out[50];

assign \d_out_out[51]~input_o  = d_out_out[51];

assign \d_out_out[52]~input_o  = d_out_out[52];

assign \d_out_out[53]~input_o  = d_out_out[53];

assign \d_out_out[54]~input_o  = d_out_out[54];

assign \d_out_out[55]~input_o  = d_out_out[55];

assign \d_out_out[56]~input_o  = d_out_out[56];

assign \d_out_out[57]~input_o  = d_out_out[57];

assign \d_out_out[58]~input_o  = d_out_out[58];

assign \d_out_out[59]~input_o  = d_out_out[59];

assign \d_out_out[60]~input_o  = d_out_out[60];

assign \d_out_out[61]~input_o  = d_out_out[61];

assign \d_out_out[62]~input_o  = d_out_out[62];

assign \d_out_out[63]~input_o  = d_out_out[63];

assign \d_out_out[64]~input_o  = d_out_out[64];

assign \d_out_out[65]~input_o  = d_out_out[65];

assign \d_out_out[66]~input_o  = d_out_out[66];

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \ram_mm_chipselect~input_o  = ram_mm_chipselect;

assign \ram_mm_write~input_o  = ram_mm_write;

assign \ram_clk_clk~input_o  = ram_clk_clk;

assign \ram_mm_clken~input_o  = ram_mm_clken;

assign \ram_mm_writedata[0]~input_o  = ram_mm_writedata[0];

assign \ram_mm_address[0]~input_o  = ram_mm_address[0];

assign \ram_mm_address[1]~input_o  = ram_mm_address[1];

assign \ram_mm_address[2]~input_o  = ram_mm_address[2];

assign \ram_mm_address[3]~input_o  = ram_mm_address[3];

assign \ram_mm_address[4]~input_o  = ram_mm_address[4];

assign \ram_mm_address[5]~input_o  = ram_mm_address[5];

assign \ram_mm_address[6]~input_o  = ram_mm_address[6];

assign \ram_mm_address[7]~input_o  = ram_mm_address[7];

assign \ram_mm_address[8]~input_o  = ram_mm_address[8];

assign \ram_mm_address[9]~input_o  = ram_mm_address[9];

assign \ram_mm_address[10]~input_o  = ram_mm_address[10];

assign \ram_mm_address[11]~input_o  = ram_mm_address[11];

assign \ram_mm_address[12]~input_o  = ram_mm_address[12];

assign \ram_mm_byteenable[0]~input_o  = ram_mm_byteenable[0];

assign \ram_mm_writedata[1]~input_o  = ram_mm_writedata[1];

assign \ram_mm_writedata[2]~input_o  = ram_mm_writedata[2];

assign \ram_mm_writedata[3]~input_o  = ram_mm_writedata[3];

assign \ram_mm_writedata[4]~input_o  = ram_mm_writedata[4];

assign \ram_mm_writedata[5]~input_o  = ram_mm_writedata[5];

assign \ram_mm_writedata[6]~input_o  = ram_mm_writedata[6];

assign \ram_mm_writedata[7]~input_o  = ram_mm_writedata[7];

assign \ram_mm_writedata[8]~input_o  = ram_mm_writedata[8];

assign \ram_mm_byteenable[1]~input_o  = ram_mm_byteenable[1];

assign \ram_mm_writedata[9]~input_o  = ram_mm_writedata[9];

assign \ram_mm_writedata[10]~input_o  = ram_mm_writedata[10];

assign \ram_mm_writedata[11]~input_o  = ram_mm_writedata[11];

assign \ram_mm_writedata[12]~input_o  = ram_mm_writedata[12];

assign \ram_mm_writedata[13]~input_o  = ram_mm_writedata[13];

assign \ram_mm_writedata[14]~input_o  = ram_mm_writedata[14];

assign \ram_mm_writedata[15]~input_o  = ram_mm_writedata[15];

assign \ram_mm_writedata[16]~input_o  = ram_mm_writedata[16];

assign \ram_mm_byteenable[2]~input_o  = ram_mm_byteenable[2];

assign \ram_mm_writedata[17]~input_o  = ram_mm_writedata[17];

assign \ram_mm_writedata[18]~input_o  = ram_mm_writedata[18];

assign \ram_mm_writedata[19]~input_o  = ram_mm_writedata[19];

assign \ram_mm_writedata[20]~input_o  = ram_mm_writedata[20];

assign \ram_mm_writedata[21]~input_o  = ram_mm_writedata[21];

assign \ram_mm_writedata[22]~input_o  = ram_mm_writedata[22];

assign \ram_mm_writedata[23]~input_o  = ram_mm_writedata[23];

assign \ram_mm_writedata[24]~input_o  = ram_mm_writedata[24];

assign \ram_mm_byteenable[3]~input_o  = ram_mm_byteenable[3];

assign \ram_mm_writedata[25]~input_o  = ram_mm_writedata[25];

assign \ram_mm_writedata[26]~input_o  = ram_mm_writedata[26];

assign \ram_mm_writedata[27]~input_o  = ram_mm_writedata[27];

assign \ram_mm_writedata[28]~input_o  = ram_mm_writedata[28];

assign \ram_mm_writedata[29]~input_o  = ram_mm_writedata[29];

assign \ram_mm_writedata[30]~input_o  = ram_mm_writedata[30];

assign \ram_mm_writedata[31]~input_o  = ram_mm_writedata[31];

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck_n),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_spim0_inst_MOSI[0]~output (
	.i(\hps_0|hps_io|border|intermediate[36] ),
	.oe(\hps_0|hps_io|border|intermediate[37] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_spim0_inst_MOSI),
	.obar());
defparam \hps_0|hps_io|border|hps_io_spim0_inst_MOSI[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_spim0_inst_MOSI[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_spim0_inst_MOSI[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output (
	.i(\hps_0|hps_io|border|intermediate[38] ),
	.oe(\hps_0|hps_io|border|intermediate[39] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_spim1_inst_MOSI),
	.obar());
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .shift_series_termination_control = "false";

assign clk_100m_clk = \pll_0|altera_pll_i|outclk_wire[0] ;

assign d_out_in[0] = \hps_0|fpga_interfaces|h2f_loan_in[0] ;

assign d_out_in[1] = \hps_0|fpga_interfaces|h2f_loan_in[1] ;

assign d_out_in[2] = \hps_0|fpga_interfaces|h2f_loan_in[2] ;

assign d_out_in[3] = \hps_0|fpga_interfaces|h2f_loan_in[3] ;

assign d_out_in[4] = \hps_0|fpga_interfaces|h2f_loan_in[4] ;

assign d_out_in[5] = \hps_0|fpga_interfaces|h2f_loan_in[5] ;

assign d_out_in[6] = \hps_0|fpga_interfaces|h2f_loan_in[6] ;

assign d_out_in[7] = \hps_0|fpga_interfaces|h2f_loan_in[7] ;

assign d_out_in[8] = \hps_0|fpga_interfaces|h2f_loan_in[8] ;

assign d_out_in[9] = \hps_0|fpga_interfaces|h2f_loan_in[9] ;

assign d_out_in[10] = \hps_0|fpga_interfaces|h2f_loan_in[10] ;

assign d_out_in[11] = \hps_0|fpga_interfaces|h2f_loan_in[11] ;

assign d_out_in[12] = \hps_0|fpga_interfaces|h2f_loan_in[12] ;

assign d_out_in[13] = \hps_0|fpga_interfaces|h2f_loan_in[13] ;

assign d_out_in[14] = \hps_0|fpga_interfaces|h2f_loan_in[14] ;

assign d_out_in[15] = \hps_0|fpga_interfaces|h2f_loan_in[15] ;

assign d_out_in[16] = \hps_0|fpga_interfaces|h2f_loan_in[16] ;

assign d_out_in[17] = \hps_0|fpga_interfaces|h2f_loan_in[17] ;

assign d_out_in[18] = \hps_0|fpga_interfaces|h2f_loan_in[18] ;

assign d_out_in[19] = \hps_0|fpga_interfaces|h2f_loan_in[19] ;

assign d_out_in[20] = \hps_0|fpga_interfaces|h2f_loan_in[20] ;

assign d_out_in[21] = \hps_0|fpga_interfaces|h2f_loan_in[21] ;

assign d_out_in[22] = \hps_0|fpga_interfaces|h2f_loan_in[22] ;

assign d_out_in[23] = \hps_0|fpga_interfaces|h2f_loan_in[23] ;

assign d_out_in[24] = \hps_0|fpga_interfaces|h2f_loan_in[24] ;

assign d_out_in[25] = \hps_0|fpga_interfaces|h2f_loan_in[25] ;

assign d_out_in[26] = \hps_0|fpga_interfaces|h2f_loan_in[26] ;

assign d_out_in[27] = \hps_0|fpga_interfaces|h2f_loan_in[27] ;

assign d_out_in[28] = \hps_0|fpga_interfaces|h2f_loan_in[28] ;

assign d_out_in[29] = \hps_0|fpga_interfaces|h2f_loan_in[29] ;

assign d_out_in[30] = \hps_0|fpga_interfaces|h2f_loan_in[30] ;

assign d_out_in[31] = \hps_0|fpga_interfaces|h2f_loan_in[31] ;

assign d_out_in[32] = \hps_0|fpga_interfaces|h2f_loan_in[32] ;

assign d_out_in[33] = \hps_0|fpga_interfaces|h2f_loan_in[33] ;

assign d_out_in[34] = \hps_0|fpga_interfaces|h2f_loan_in[34] ;

assign d_out_in[35] = \hps_0|fpga_interfaces|h2f_loan_in[35] ;

assign d_out_in[36] = \hps_0|fpga_interfaces|h2f_loan_in[36] ;

assign d_out_in[37] = \hps_0|fpga_interfaces|h2f_loan_in[37] ;

assign d_out_in[38] = \hps_0|fpga_interfaces|h2f_loan_in[38] ;

assign d_out_in[39] = \hps_0|fpga_interfaces|h2f_loan_in[39] ;

assign d_out_in[40] = \hps_0|fpga_interfaces|h2f_loan_in[40] ;

assign d_out_in[41] = \hps_0|fpga_interfaces|h2f_loan_in[41] ;

assign d_out_in[42] = \hps_0|fpga_interfaces|h2f_loan_in[42] ;

assign d_out_in[43] = \hps_0|fpga_interfaces|h2f_loan_in[43] ;

assign d_out_in[44] = \hps_0|fpga_interfaces|h2f_loan_in[44] ;

assign d_out_in[45] = \hps_0|fpga_interfaces|h2f_loan_in[45] ;

assign d_out_in[46] = \hps_0|fpga_interfaces|h2f_loan_in[46] ;

assign d_out_in[47] = \hps_0|fpga_interfaces|h2f_loan_in[47] ;

assign d_out_in[48] = \hps_0|fpga_interfaces|h2f_loan_in[48] ;

assign d_out_in[49] = \hps_0|fpga_interfaces|h2f_loan_in[49] ;

assign d_out_in[50] = \hps_0|fpga_interfaces|h2f_loan_in[50] ;

assign d_out_in[51] = \hps_0|fpga_interfaces|h2f_loan_in[51] ;

assign d_out_in[52] = \hps_0|fpga_interfaces|h2f_loan_in[52] ;

assign d_out_in[53] = \hps_0|fpga_interfaces|h2f_loan_in[53] ;

assign d_out_in[54] = \hps_0|fpga_interfaces|h2f_loan_in[54] ;

assign d_out_in[55] = \hps_0|fpga_interfaces|h2f_loan_in[55] ;

assign d_out_in[56] = \hps_0|fpga_interfaces|h2f_loan_in[56] ;

assign d_out_in[57] = \hps_0|fpga_interfaces|h2f_loan_in[57] ;

assign d_out_in[58] = \hps_0|fpga_interfaces|h2f_loan_in[58] ;

assign d_out_in[59] = \hps_0|fpga_interfaces|h2f_loan_in[59] ;

assign d_out_in[60] = \hps_0|fpga_interfaces|h2f_loan_in[60] ;

assign d_out_in[61] = \hps_0|fpga_interfaces|h2f_loan_in[61] ;

assign d_out_in[62] = \hps_0|fpga_interfaces|h2f_loan_in[62] ;

assign d_out_in[63] = \hps_0|fpga_interfaces|h2f_loan_in[63] ;

assign d_out_in[64] = \hps_0|fpga_interfaces|h2f_loan_in[64] ;

assign d_out_in[65] = \hps_0|fpga_interfaces|h2f_loan_in[65] ;

assign d_out_in[66] = \hps_0|fpga_interfaces|h2f_loan_in[66] ;

assign hps_io_hps_io_emac1_inst_TX_CLK = \hps_0|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;

assign hps_io_hps_io_emac1_inst_TXD0 = \hps_0|hps_io|border|emac1_inst~emac_phy_txd ;

assign hps_io_hps_io_emac1_inst_TXD1 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;

assign hps_io_hps_io_emac1_inst_TXD2 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;

assign hps_io_hps_io_emac1_inst_TXD3 = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;

assign hps_io_hps_io_emac1_inst_MDC = \hps_0|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;

assign hps_io_hps_io_emac1_inst_TX_CTL = \hps_0|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;

assign hps_io_hps_io_qspi_inst_SS0 = \hps_0|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;

assign hps_io_hps_io_qspi_inst_CLK = \hps_0|hps_io|border|qspi_inst~O_QSPI_SCLK ;

assign hps_io_hps_io_sdio_inst_CLK = \hps_0|hps_io|border|sdio_inst~sdmmc_cclk ;

assign hps_io_hps_io_usb1_inst_STP = \hps_0|hps_io|border|usb1_inst~usb_ulpi_stp ;

assign hps_io_hps_io_spim0_inst_CLK = \hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SCLK ;

assign hps_io_hps_io_spim0_inst_SS0 = \hps_0|hps_io|border|spim0_inst~O_SPI_MASTER_SS_0_N ;

assign hps_io_hps_io_spim1_inst_CLK = \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;

assign hps_io_hps_io_spim1_inst_SS0 = \hps_0|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;

assign hps_io_hps_io_uart0_inst_TX = \hps_0|hps_io|border|uart0_inst~uart_txd ;

assign memory_mem_a[0] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;

assign memory_mem_a[1] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;

assign memory_mem_a[2] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;

assign memory_mem_a[3] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;

assign memory_mem_a[4] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;

assign memory_mem_a[5] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;

assign memory_mem_a[6] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;

assign memory_mem_a[7] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;

assign memory_mem_a[8] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;

assign memory_mem_a[9] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;

assign memory_mem_a[10] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;

assign memory_mem_a[11] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;

assign memory_mem_a[12] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;

assign memory_mem_a[13] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;

assign memory_mem_a[14] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;

assign memory_mem_ba[0] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;

assign memory_mem_ba[1] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;

assign memory_mem_ba[2] = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;

assign memory_mem_cke = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;

assign memory_mem_cs_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;

assign memory_mem_ras_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;

assign memory_mem_cas_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;

assign memory_mem_we_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;

assign memory_mem_reset_n = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;

assign memory_mem_odt = \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;

assign ram_mm_readdata[0] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[0] ;

assign ram_mm_readdata[1] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[1] ;

assign ram_mm_readdata[2] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[2] ;

assign ram_mm_readdata[3] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[3] ;

assign ram_mm_readdata[4] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[4] ;

assign ram_mm_readdata[5] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[5] ;

assign ram_mm_readdata[6] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[6] ;

assign ram_mm_readdata[7] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[7] ;

assign ram_mm_readdata[8] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[8] ;

assign ram_mm_readdata[9] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[9] ;

assign ram_mm_readdata[10] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[10] ;

assign ram_mm_readdata[11] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[11] ;

assign ram_mm_readdata[12] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[12] ;

assign ram_mm_readdata[13] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[13] ;

assign ram_mm_readdata[14] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[14] ;

assign ram_mm_readdata[15] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[15] ;

assign ram_mm_readdata[16] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[16] ;

assign ram_mm_readdata[17] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[17] ;

assign ram_mm_readdata[18] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[18] ;

assign ram_mm_readdata[19] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[19] ;

assign ram_mm_readdata[20] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[20] ;

assign ram_mm_readdata[21] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[21] ;

assign ram_mm_readdata[22] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[22] ;

assign ram_mm_readdata[23] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[23] ;

assign ram_mm_readdata[24] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[24] ;

assign ram_mm_readdata[25] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[25] ;

assign ram_mm_readdata[26] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[26] ;

assign ram_mm_readdata[27] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[27] ;

assign ram_mm_readdata[28] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[28] ;

assign ram_mm_readdata[29] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[29] ;

assign ram_mm_readdata[30] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[30] ;

assign ram_mm_readdata[31] = \onchip_memory2_0|the_altsyncram|auto_generated|q_b[31] ;

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output (
	.i(\hps_0|hps_io|border|intermediate[0] ),
	.oe(\hps_0|hps_io|border|intermediate[1] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_emac1_inst_MDIO),
	.obar());
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[2] ),
	.oe(\hps_0|hps_io|border|intermediate[3] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[4] ),
	.oe(\hps_0|hps_io|border|intermediate[5] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[6] ),
	.oe(\hps_0|hps_io|border|intermediate[7] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[8] ),
	.oe(\hps_0|hps_io|border|intermediate[9] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_qspi_inst_IO3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output (
	.i(\hps_0|hps_io|border|intermediate[10] ),
	.oe(\hps_0|hps_io|border|intermediate[11] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_CMD),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_CMD[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[12] ),
	.oe(\hps_0|hps_io|border|intermediate[13] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[14] ),
	.oe(\hps_0|hps_io|border|intermediate[15] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[16] ),
	.oe(\hps_0|hps_io|border|intermediate[17] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[18] ),
	.oe(\hps_0|hps_io|border|intermediate[19] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_sdio_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output (
	.i(\hps_0|hps_io|border|intermediate[20] ),
	.oe(\hps_0|hps_io|border|intermediate[21] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D0),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output (
	.i(\hps_0|hps_io|border|intermediate[22] ),
	.oe(\hps_0|hps_io|border|intermediate[23] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D1),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output (
	.i(\hps_0|hps_io|border|intermediate[24] ),
	.oe(\hps_0|hps_io|border|intermediate[25] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D2),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output (
	.i(\hps_0|hps_io|border|intermediate[26] ),
	.oe(\hps_0|hps_io|border|intermediate[27] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D3),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output (
	.i(\hps_0|hps_io|border|intermediate[28] ),
	.oe(\hps_0|hps_io|border|intermediate[29] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D4),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D4[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output (
	.i(\hps_0|hps_io|border|intermediate[30] ),
	.oe(\hps_0|hps_io|border|intermediate[31] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D5),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D5[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output (
	.i(\hps_0|hps_io|border|intermediate[32] ),
	.oe(\hps_0|hps_io|border|intermediate[33] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D6),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D6[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output (
	.i(\hps_0|hps_io|border|intermediate[34] ),
	.oe(\hps_0|hps_io|border|intermediate[35] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D7),
	.obar());
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_usb1_inst_D7[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output (
	.i(\hps_0|hps_io|border|intermediate[40] ),
	.oe(\hps_0|hps_io|border|intermediate[41] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO09),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output (
	.i(\hps_0|hps_io|border|intermediate[42] ),
	.oe(\hps_0|hps_io|border|intermediate[43] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO40),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output (
	.i(\hps_0|hps_io|border|intermediate[44] ),
	.oe(\hps_0|hps_io|border|intermediate[45] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO48),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output (
	.i(\hps_0|hps_io|border|intermediate[46] ),
	.oe(\hps_0|hps_io|border|intermediate[47] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO61),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~output (
	.i(\hps_0|hps_io|border|intermediate[48] ),
	.oe(\hps_0|hps_io|border|intermediate[49] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO62),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_GPIO62[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~output (
	.i(\hps_0|hps_io|border|intermediate[50] ),
	.oe(\hps_0|hps_io|border|intermediate[51] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO00),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO00[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~output (
	.i(\hps_0|hps_io|border|intermediate[52] ),
	.oe(\hps_0|hps_io|border|intermediate[53] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO41),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO41[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~output (
	.i(\hps_0|hps_io|border|intermediate[54] ),
	.oe(\hps_0|hps_io|border|intermediate[55] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO51),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO51[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~output (
	.i(\hps_0|hps_io|border|intermediate[56] ),
	.oe(\hps_0|hps_io|border|intermediate[57] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO52),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO52[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~output (
	.i(\hps_0|hps_io|border|intermediate[58] ),
	.oe(\hps_0|hps_io|border|intermediate[59] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO53),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO53[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~output (
	.i(\hps_0|hps_io|border|intermediate[60] ),
	.oe(\hps_0|hps_io|border|intermediate[61] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO54),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO54[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~output (
	.i(\hps_0|hps_io|border|intermediate[62] ),
	.oe(\hps_0|hps_io|border|intermediate[63] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO55),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO55[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~output (
	.i(\hps_0|hps_io|border|intermediate[64] ),
	.oe(\hps_0|hps_io|border|intermediate[65] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_LOANIO56),
	.obar());
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~output .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~output .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_io_gpio_inst_LOANIO56[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[4]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[5]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[6]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[7]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[8]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[9]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[10]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[11]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[12]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[13]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[14]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[15]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[16]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[17]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[18]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[19]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[20]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[21]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[22]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[23]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[24]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[25]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[26]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[27]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[28]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[29]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[30]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[31]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[0]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[1]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[2]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps_0|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[3]),
	.obar());
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps_0|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

assign \ram_reset_reset~input_o  = ram_reset_reset;

endmodule

module soc_system_altera_reset_controller (
	outclk_wire_0,
	altera_reset_synchronizer_int_chain_out,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.reset_reset_n(reset_reset_n));

endmodule

module soc_system_altera_reset_controller_1 (
	h2f_rst_n_0,
	outclk_wire_0,
	altera_reset_synchronizer_int_chain_out)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	outclk_wire_0;
output 	altera_reset_synchronizer_int_chain_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out));

endmodule

module soc_system_altera_reset_synchronizer_1 (
	h2f_rst_n_0,
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module soc_system_altera_reset_synchronizer_3 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module soc_system_soc_system_hps_0 (
	h2f_loan_in_0,
	h2f_loan_in_1,
	h2f_loan_in_2,
	h2f_loan_in_3,
	h2f_loan_in_4,
	h2f_loan_in_5,
	h2f_loan_in_6,
	h2f_loan_in_7,
	h2f_loan_in_8,
	h2f_loan_in_9,
	h2f_loan_in_10,
	h2f_loan_in_11,
	h2f_loan_in_12,
	h2f_loan_in_13,
	h2f_loan_in_14,
	h2f_loan_in_15,
	h2f_loan_in_16,
	h2f_loan_in_17,
	h2f_loan_in_18,
	h2f_loan_in_19,
	h2f_loan_in_20,
	h2f_loan_in_21,
	h2f_loan_in_22,
	h2f_loan_in_23,
	h2f_loan_in_24,
	h2f_loan_in_25,
	h2f_loan_in_26,
	h2f_loan_in_27,
	h2f_loan_in_28,
	h2f_loan_in_29,
	h2f_loan_in_30,
	h2f_loan_in_31,
	h2f_loan_in_32,
	h2f_loan_in_33,
	h2f_loan_in_34,
	h2f_loan_in_35,
	h2f_loan_in_36,
	h2f_loan_in_37,
	h2f_loan_in_38,
	h2f_loan_in_39,
	h2f_loan_in_40,
	h2f_loan_in_41,
	h2f_loan_in_42,
	h2f_loan_in_43,
	h2f_loan_in_44,
	h2f_loan_in_45,
	h2f_loan_in_46,
	h2f_loan_in_47,
	h2f_loan_in_48,
	h2f_loan_in_49,
	h2f_loan_in_50,
	h2f_loan_in_51,
	h2f_loan_in_52,
	h2f_loan_in_53,
	h2f_loan_in_54,
	h2f_loan_in_55,
	h2f_loan_in_56,
	h2f_loan_in_57,
	h2f_loan_in_58,
	h2f_loan_in_59,
	h2f_loan_in_60,
	h2f_loan_in_61,
	h2f_loan_in_62,
	h2f_loan_in_63,
	h2f_loan_in_64,
	h2f_loan_in_65,
	h2f_loan_in_66,
	h2f_rst_n_0,
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	sink1_ready,
	awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	wready,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim0_inst,
	spim0_inst1,
	intermediate_36,
	intermediate_37,
	spim1_inst,
	spim1_inst1,
	intermediate_38,
	intermediate_39,
	uart0_inst,
	intermediate_50,
	intermediate_40,
	intermediate_51,
	intermediate_41,
	intermediate_42,
	intermediate_52,
	intermediate_44,
	intermediate_54,
	intermediate_56,
	intermediate_58,
	intermediate_60,
	intermediate_62,
	intermediate_64,
	intermediate_43,
	intermediate_53,
	intermediate_45,
	intermediate_55,
	intermediate_57,
	intermediate_59,
	intermediate_61,
	intermediate_63,
	intermediate_65,
	intermediate_46,
	intermediate_48,
	intermediate_47,
	intermediate_49,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_gpio_inst_GPIO62_0,
	hps_io_gpio_inst_LOANIO00_0,
	hps_io_gpio_inst_LOANIO41_0,
	hps_io_gpio_inst_LOANIO51_0,
	hps_io_gpio_inst_LOANIO52_0,
	hps_io_gpio_inst_LOANIO53_0,
	hps_io_gpio_inst_LOANIO54_0,
	hps_io_gpio_inst_LOANIO55_0,
	hps_io_gpio_inst_LOANIO56_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim0_inst_MISO,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin,
	d_out_oe_0,
	d_out_oe_1,
	d_out_oe_2,
	d_out_oe_3,
	d_out_oe_4,
	d_out_oe_5,
	d_out_oe_6,
	d_out_oe_7,
	d_out_oe_8,
	d_out_oe_9,
	d_out_oe_10,
	d_out_oe_11,
	d_out_oe_12,
	d_out_oe_13,
	d_out_oe_14,
	d_out_oe_15,
	d_out_oe_16,
	d_out_oe_17,
	d_out_oe_18,
	d_out_oe_19,
	d_out_oe_20,
	d_out_oe_21,
	d_out_oe_22,
	d_out_oe_23,
	d_out_oe_24,
	d_out_oe_25,
	d_out_oe_26,
	d_out_oe_27,
	d_out_oe_28,
	d_out_oe_29,
	d_out_oe_30,
	d_out_oe_31,
	d_out_oe_32,
	d_out_oe_33,
	d_out_oe_34,
	d_out_oe_35,
	d_out_oe_36,
	d_out_oe_37,
	d_out_oe_38,
	d_out_oe_39,
	d_out_oe_40,
	d_out_oe_41,
	d_out_oe_42,
	d_out_oe_43,
	d_out_oe_44,
	d_out_oe_45,
	d_out_oe_46,
	d_out_oe_47,
	d_out_oe_48,
	d_out_oe_49,
	d_out_oe_50,
	d_out_oe_51,
	d_out_oe_52,
	d_out_oe_53,
	d_out_oe_54,
	d_out_oe_55,
	d_out_oe_56,
	d_out_oe_57,
	d_out_oe_58,
	d_out_oe_59,
	d_out_oe_60,
	d_out_oe_61,
	d_out_oe_62,
	d_out_oe_63,
	d_out_oe_64,
	d_out_oe_65,
	d_out_oe_66,
	d_out_out_0,
	d_out_out_1,
	d_out_out_2,
	d_out_out_3,
	d_out_out_4,
	d_out_out_5,
	d_out_out_6,
	d_out_out_7,
	d_out_out_8,
	d_out_out_9,
	d_out_out_10,
	d_out_out_11,
	d_out_out_12,
	d_out_out_13,
	d_out_out_14,
	d_out_out_15,
	d_out_out_16,
	d_out_out_17,
	d_out_out_18,
	d_out_out_19,
	d_out_out_20,
	d_out_out_21,
	d_out_out_22,
	d_out_out_23,
	d_out_out_24,
	d_out_out_25,
	d_out_out_26,
	d_out_out_27,
	d_out_out_28,
	d_out_out_29,
	d_out_out_30,
	d_out_out_31,
	d_out_out_32,
	d_out_out_33,
	d_out_out_34,
	d_out_out_35,
	d_out_out_36,
	d_out_out_37,
	d_out_out_38,
	d_out_out_39,
	d_out_out_40,
	d_out_out_41,
	d_out_out_42,
	d_out_out_43,
	d_out_out_44,
	d_out_out_45,
	d_out_out_46,
	d_out_out_47,
	d_out_out_48,
	d_out_out_49,
	d_out_out_50,
	d_out_out_51,
	d_out_out_52,
	d_out_out_53,
	d_out_out_54,
	d_out_out_55,
	d_out_out_56,
	d_out_out_57,
	d_out_out_58,
	d_out_out_59,
	d_out_out_60,
	d_out_out_61,
	d_out_out_62,
	d_out_out_63,
	d_out_out_64,
	d_out_out_65,
	d_out_out_66)/* synthesis synthesis_greybox=0 */;
output 	h2f_loan_in_0;
output 	h2f_loan_in_1;
output 	h2f_loan_in_2;
output 	h2f_loan_in_3;
output 	h2f_loan_in_4;
output 	h2f_loan_in_5;
output 	h2f_loan_in_6;
output 	h2f_loan_in_7;
output 	h2f_loan_in_8;
output 	h2f_loan_in_9;
output 	h2f_loan_in_10;
output 	h2f_loan_in_11;
output 	h2f_loan_in_12;
output 	h2f_loan_in_13;
output 	h2f_loan_in_14;
output 	h2f_loan_in_15;
output 	h2f_loan_in_16;
output 	h2f_loan_in_17;
output 	h2f_loan_in_18;
output 	h2f_loan_in_19;
output 	h2f_loan_in_20;
output 	h2f_loan_in_21;
output 	h2f_loan_in_22;
output 	h2f_loan_in_23;
output 	h2f_loan_in_24;
output 	h2f_loan_in_25;
output 	h2f_loan_in_26;
output 	h2f_loan_in_27;
output 	h2f_loan_in_28;
output 	h2f_loan_in_29;
output 	h2f_loan_in_30;
output 	h2f_loan_in_31;
output 	h2f_loan_in_32;
output 	h2f_loan_in_33;
output 	h2f_loan_in_34;
output 	h2f_loan_in_35;
output 	h2f_loan_in_36;
output 	h2f_loan_in_37;
output 	h2f_loan_in_38;
output 	h2f_loan_in_39;
output 	h2f_loan_in_40;
output 	h2f_loan_in_41;
output 	h2f_loan_in_42;
output 	h2f_loan_in_43;
output 	h2f_loan_in_44;
output 	h2f_loan_in_45;
output 	h2f_loan_in_46;
output 	h2f_loan_in_47;
output 	h2f_loan_in_48;
output 	h2f_loan_in_49;
output 	h2f_loan_in_50;
output 	h2f_loan_in_51;
output 	h2f_loan_in_52;
output 	h2f_loan_in_53;
output 	h2f_loan_in_54;
output 	h2f_loan_in_55;
output 	h2f_loan_in_56;
output 	h2f_loan_in_57;
output 	h2f_loan_in_58;
output 	h2f_loan_in_59;
output 	h2f_loan_in_60;
output 	h2f_loan_in_61;
output 	h2f_loan_in_62;
output 	h2f_loan_in_63;
output 	h2f_loan_in_64;
output 	h2f_loan_in_65;
output 	h2f_loan_in_66;
output 	h2f_rst_n_0;
output 	h2f_lw_ARVALID_0;
output 	h2f_lw_AWVALID_0;
output 	h2f_lw_BREADY_0;
output 	h2f_lw_RREADY_0;
output 	h2f_lw_WLAST_0;
output 	h2f_lw_WVALID_0;
output 	h2f_lw_ARADDR_0;
output 	h2f_lw_ARADDR_1;
output 	h2f_lw_ARADDR_2;
output 	h2f_lw_ARADDR_3;
output 	h2f_lw_ARADDR_4;
output 	h2f_lw_ARADDR_5;
output 	h2f_lw_ARADDR_6;
output 	h2f_lw_ARADDR_7;
output 	h2f_lw_ARADDR_8;
output 	h2f_lw_ARADDR_9;
output 	h2f_lw_ARADDR_10;
output 	h2f_lw_ARADDR_11;
output 	h2f_lw_ARADDR_12;
output 	h2f_lw_ARADDR_13;
output 	h2f_lw_ARADDR_14;
output 	h2f_lw_ARBURST_0;
output 	h2f_lw_ARBURST_1;
output 	h2f_lw_ARID_0;
output 	h2f_lw_ARID_1;
output 	h2f_lw_ARID_2;
output 	h2f_lw_ARID_3;
output 	h2f_lw_ARID_4;
output 	h2f_lw_ARID_5;
output 	h2f_lw_ARID_6;
output 	h2f_lw_ARID_7;
output 	h2f_lw_ARID_8;
output 	h2f_lw_ARID_9;
output 	h2f_lw_ARID_10;
output 	h2f_lw_ARID_11;
output 	h2f_lw_ARLEN_0;
output 	h2f_lw_ARLEN_1;
output 	h2f_lw_ARLEN_2;
output 	h2f_lw_ARLEN_3;
output 	h2f_lw_ARSIZE_0;
output 	h2f_lw_ARSIZE_1;
output 	h2f_lw_ARSIZE_2;
output 	h2f_lw_AWADDR_0;
output 	h2f_lw_AWADDR_1;
output 	h2f_lw_AWADDR_2;
output 	h2f_lw_AWADDR_3;
output 	h2f_lw_AWADDR_4;
output 	h2f_lw_AWADDR_5;
output 	h2f_lw_AWADDR_6;
output 	h2f_lw_AWADDR_7;
output 	h2f_lw_AWADDR_8;
output 	h2f_lw_AWADDR_9;
output 	h2f_lw_AWADDR_10;
output 	h2f_lw_AWADDR_11;
output 	h2f_lw_AWADDR_12;
output 	h2f_lw_AWADDR_13;
output 	h2f_lw_AWADDR_14;
output 	h2f_lw_AWBURST_0;
output 	h2f_lw_AWBURST_1;
output 	h2f_lw_AWID_0;
output 	h2f_lw_AWID_1;
output 	h2f_lw_AWID_2;
output 	h2f_lw_AWID_3;
output 	h2f_lw_AWID_4;
output 	h2f_lw_AWID_5;
output 	h2f_lw_AWID_6;
output 	h2f_lw_AWID_7;
output 	h2f_lw_AWID_8;
output 	h2f_lw_AWID_9;
output 	h2f_lw_AWID_10;
output 	h2f_lw_AWID_11;
output 	h2f_lw_AWLEN_0;
output 	h2f_lw_AWLEN_1;
output 	h2f_lw_AWLEN_2;
output 	h2f_lw_AWLEN_3;
output 	h2f_lw_AWSIZE_0;
output 	h2f_lw_AWSIZE_1;
output 	h2f_lw_AWSIZE_2;
output 	h2f_lw_WDATA_0;
output 	h2f_lw_WDATA_1;
output 	h2f_lw_WDATA_2;
output 	h2f_lw_WDATA_3;
output 	h2f_lw_WDATA_4;
output 	h2f_lw_WDATA_5;
output 	h2f_lw_WDATA_6;
output 	h2f_lw_WDATA_7;
output 	h2f_lw_WDATA_8;
output 	h2f_lw_WDATA_9;
output 	h2f_lw_WDATA_10;
output 	h2f_lw_WDATA_11;
output 	h2f_lw_WDATA_12;
output 	h2f_lw_WDATA_13;
output 	h2f_lw_WDATA_14;
output 	h2f_lw_WDATA_15;
output 	h2f_lw_WDATA_16;
output 	h2f_lw_WDATA_17;
output 	h2f_lw_WDATA_18;
output 	h2f_lw_WDATA_19;
output 	h2f_lw_WDATA_20;
output 	h2f_lw_WDATA_21;
output 	h2f_lw_WDATA_22;
output 	h2f_lw_WDATA_23;
output 	h2f_lw_WDATA_24;
output 	h2f_lw_WDATA_25;
output 	h2f_lw_WDATA_26;
output 	h2f_lw_WDATA_27;
output 	h2f_lw_WDATA_28;
output 	h2f_lw_WDATA_29;
output 	h2f_lw_WDATA_30;
output 	h2f_lw_WDATA_31;
output 	h2f_lw_WSTRB_0;
output 	h2f_lw_WSTRB_1;
output 	h2f_lw_WSTRB_2;
output 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	sink1_ready;
input 	awready;
input 	src0_valid;
input 	source_endofpacket;
input 	src1_valid;
input 	wready;
input 	mem_88_0;
input 	mem_89_0;
input 	mem_90_0;
input 	mem_91_0;
input 	mem_92_0;
input 	mem_93_0;
input 	mem_94_0;
input 	mem_95_0;
input 	mem_96_0;
input 	mem_97_0;
input 	mem_98_0;
input 	mem_99_0;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	out_data_8;
input 	out_data_9;
input 	out_data_10;
input 	out_data_11;
input 	out_data_12;
input 	out_data_13;
input 	out_data_14;
input 	out_data_15;
input 	out_data_16;
input 	out_data_17;
input 	out_data_18;
input 	out_data_19;
input 	out_data_20;
input 	out_data_21;
input 	out_data_22;
input 	out_data_23;
input 	out_data_24;
input 	out_data_25;
input 	out_data_26;
input 	out_data_27;
input 	out_data_28;
input 	out_data_29;
input 	out_data_30;
input 	out_data_31;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim0_inst;
output 	spim0_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_38;
output 	intermediate_39;
output 	uart0_inst;
output 	intermediate_50;
output 	intermediate_40;
output 	intermediate_51;
output 	intermediate_41;
output 	intermediate_42;
output 	intermediate_52;
output 	intermediate_44;
output 	intermediate_54;
output 	intermediate_56;
output 	intermediate_58;
output 	intermediate_60;
output 	intermediate_62;
output 	intermediate_64;
output 	intermediate_43;
output 	intermediate_53;
output 	intermediate_45;
output 	intermediate_55;
output 	intermediate_57;
output 	intermediate_59;
output 	intermediate_61;
output 	intermediate_63;
output 	intermediate_65;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_47;
output 	intermediate_49;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_gpio_inst_GPIO62_0;
input 	hps_io_gpio_inst_LOANIO00_0;
input 	hps_io_gpio_inst_LOANIO41_0;
input 	hps_io_gpio_inst_LOANIO51_0;
input 	hps_io_gpio_inst_LOANIO52_0;
input 	hps_io_gpio_inst_LOANIO53_0;
input 	hps_io_gpio_inst_LOANIO54_0;
input 	hps_io_gpio_inst_LOANIO55_0;
input 	hps_io_gpio_inst_LOANIO56_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim0_inst_MISO;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;
input 	d_out_oe_0;
input 	d_out_oe_1;
input 	d_out_oe_2;
input 	d_out_oe_3;
input 	d_out_oe_4;
input 	d_out_oe_5;
input 	d_out_oe_6;
input 	d_out_oe_7;
input 	d_out_oe_8;
input 	d_out_oe_9;
input 	d_out_oe_10;
input 	d_out_oe_11;
input 	d_out_oe_12;
input 	d_out_oe_13;
input 	d_out_oe_14;
input 	d_out_oe_15;
input 	d_out_oe_16;
input 	d_out_oe_17;
input 	d_out_oe_18;
input 	d_out_oe_19;
input 	d_out_oe_20;
input 	d_out_oe_21;
input 	d_out_oe_22;
input 	d_out_oe_23;
input 	d_out_oe_24;
input 	d_out_oe_25;
input 	d_out_oe_26;
input 	d_out_oe_27;
input 	d_out_oe_28;
input 	d_out_oe_29;
input 	d_out_oe_30;
input 	d_out_oe_31;
input 	d_out_oe_32;
input 	d_out_oe_33;
input 	d_out_oe_34;
input 	d_out_oe_35;
input 	d_out_oe_36;
input 	d_out_oe_37;
input 	d_out_oe_38;
input 	d_out_oe_39;
input 	d_out_oe_40;
input 	d_out_oe_41;
input 	d_out_oe_42;
input 	d_out_oe_43;
input 	d_out_oe_44;
input 	d_out_oe_45;
input 	d_out_oe_46;
input 	d_out_oe_47;
input 	d_out_oe_48;
input 	d_out_oe_49;
input 	d_out_oe_50;
input 	d_out_oe_51;
input 	d_out_oe_52;
input 	d_out_oe_53;
input 	d_out_oe_54;
input 	d_out_oe_55;
input 	d_out_oe_56;
input 	d_out_oe_57;
input 	d_out_oe_58;
input 	d_out_oe_59;
input 	d_out_oe_60;
input 	d_out_oe_61;
input 	d_out_oe_62;
input 	d_out_oe_63;
input 	d_out_oe_64;
input 	d_out_oe_65;
input 	d_out_oe_66;
input 	d_out_out_0;
input 	d_out_out_1;
input 	d_out_out_2;
input 	d_out_out_3;
input 	d_out_out_4;
input 	d_out_out_5;
input 	d_out_out_6;
input 	d_out_out_7;
input 	d_out_out_8;
input 	d_out_out_9;
input 	d_out_out_10;
input 	d_out_out_11;
input 	d_out_out_12;
input 	d_out_out_13;
input 	d_out_out_14;
input 	d_out_out_15;
input 	d_out_out_16;
input 	d_out_out_17;
input 	d_out_out_18;
input 	d_out_out_19;
input 	d_out_out_20;
input 	d_out_out_21;
input 	d_out_out_22;
input 	d_out_out_23;
input 	d_out_out_24;
input 	d_out_out_25;
input 	d_out_out_26;
input 	d_out_out_27;
input 	d_out_out_28;
input 	d_out_out_29;
input 	d_out_out_30;
input 	d_out_out_31;
input 	d_out_out_32;
input 	d_out_out_33;
input 	d_out_out_34;
input 	d_out_out_35;
input 	d_out_out_36;
input 	d_out_out_37;
input 	d_out_out_38;
input 	d_out_out_39;
input 	d_out_out_40;
input 	d_out_out_41;
input 	d_out_out_42;
input 	d_out_out_43;
input 	d_out_out_44;
input 	d_out_out_45;
input 	d_out_out_46;
input 	d_out_out_47;
input 	d_out_out_48;
input 	d_out_out_49;
input 	d_out_out_50;
input 	d_out_out_51;
input 	d_out_out_52;
input 	d_out_out_53;
input 	d_out_out_54;
input 	d_out_out_55;
input 	d_out_out_56;
input 	d_out_out_57;
input 	d_out_out_58;
input 	d_out_out_59;
input 	d_out_out_60;
input 	d_out_out_61;
input 	d_out_out_62;
input 	d_out_out_63;
input 	d_out_out_64;
input 	d_out_out_65;
input 	d_out_out_66;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fpga_interfaces|loanio_gpio_loanio0_oe[0] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[1] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[2] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[3] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[4] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[5] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[6] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[7] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[8] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[9] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[10] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[11] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[12] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[13] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[14] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[15] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[16] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[17] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[18] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[19] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[20] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[21] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[22] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[23] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[24] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[25] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[26] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[27] ;
wire \fpga_interfaces|loanio_gpio_loanio0_oe[28] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[0] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[1] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[2] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[3] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[4] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[5] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[6] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[7] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[8] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[9] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[10] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[11] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[12] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[13] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[14] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[15] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[16] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[17] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[18] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[19] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[20] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[21] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[22] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[23] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[24] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[25] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[26] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[27] ;
wire \fpga_interfaces|loanio_gpio_loanio1_oe[28] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[0] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[1] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[2] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[3] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[4] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[5] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[6] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[7] ;
wire \fpga_interfaces|loanio_gpio_loanio2_oe[8] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[0] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[1] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[2] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[3] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[4] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[5] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[6] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[7] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[8] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[9] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[10] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[11] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[12] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[13] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[14] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[15] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[16] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[17] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[18] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[19] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[20] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[21] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[22] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[23] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[24] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[25] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[26] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[27] ;
wire \fpga_interfaces|loanio_gpio_loanio0_o[28] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[0] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[1] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[2] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[3] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[4] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[5] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[6] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[7] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[8] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[9] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[10] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[11] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[12] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[13] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[14] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[15] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[16] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[17] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[18] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[19] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[20] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[21] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[22] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[23] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[24] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[25] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[26] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[27] ;
wire \fpga_interfaces|loanio_gpio_loanio1_o[28] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[0] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[1] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[2] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[3] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[4] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[5] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[6] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[7] ;
wire \fpga_interfaces|loanio_gpio_loanio2_o[8] ;
wire \hps_io|border|gpio_inst~LOANIO0_I0 ;
wire \hps_io|border|gpio_inst~LOANIO0_I1 ;
wire \hps_io|border|gpio_inst~LOANIO0_I2 ;
wire \hps_io|border|gpio_inst~LOANIO0_I3 ;
wire \hps_io|border|gpio_inst~LOANIO0_I4 ;
wire \hps_io|border|gpio_inst~LOANIO0_I5 ;
wire \hps_io|border|gpio_inst~LOANIO0_I6 ;
wire \hps_io|border|gpio_inst~LOANIO0_I7 ;
wire \hps_io|border|gpio_inst~LOANIO0_I8 ;
wire \hps_io|border|gpio_inst~LOANIO0_I9 ;
wire \hps_io|border|gpio_inst~LOANIO0_I10 ;
wire \hps_io|border|gpio_inst~LOANIO0_I11 ;
wire \hps_io|border|gpio_inst~LOANIO0_I12 ;
wire \hps_io|border|gpio_inst~LOANIO0_I13 ;
wire \hps_io|border|gpio_inst~LOANIO0_I14 ;
wire \hps_io|border|gpio_inst~LOANIO0_I15 ;
wire \hps_io|border|gpio_inst~LOANIO0_I16 ;
wire \hps_io|border|gpio_inst~LOANIO0_I17 ;
wire \hps_io|border|gpio_inst~LOANIO0_I18 ;
wire \hps_io|border|gpio_inst~LOANIO0_I19 ;
wire \hps_io|border|gpio_inst~LOANIO0_I20 ;
wire \hps_io|border|gpio_inst~LOANIO0_I21 ;
wire \hps_io|border|gpio_inst~LOANIO0_I22 ;
wire \hps_io|border|gpio_inst~LOANIO0_I23 ;
wire \hps_io|border|gpio_inst~LOANIO0_I24 ;
wire \hps_io|border|gpio_inst~LOANIO0_I25 ;
wire \hps_io|border|gpio_inst~LOANIO0_I26 ;
wire \hps_io|border|gpio_inst~LOANIO0_I27 ;
wire \hps_io|border|gpio_inst~LOANIO0_I28 ;
wire \hps_io|border|gpio_inst~LOANIO1_I0 ;
wire \hps_io|border|gpio_inst~LOANIO1_I1 ;
wire \hps_io|border|gpio_inst~LOANIO1_I2 ;
wire \hps_io|border|gpio_inst~LOANIO1_I3 ;
wire \hps_io|border|gpio_inst~LOANIO1_I4 ;
wire \hps_io|border|gpio_inst~LOANIO1_I5 ;
wire \hps_io|border|gpio_inst~LOANIO1_I6 ;
wire \hps_io|border|gpio_inst~LOANIO1_I7 ;
wire \hps_io|border|gpio_inst~LOANIO1_I8 ;
wire \hps_io|border|gpio_inst~LOANIO1_I9 ;
wire \hps_io|border|gpio_inst~LOANIO1_I10 ;
wire \hps_io|border|gpio_inst~LOANIO1_I11 ;
wire \hps_io|border|gpio_inst~LOANIO1_I12 ;
wire \hps_io|border|gpio_inst~LOANIO1_I13 ;
wire \hps_io|border|gpio_inst~LOANIO1_I14 ;
wire \hps_io|border|gpio_inst~LOANIO1_I15 ;
wire \hps_io|border|gpio_inst~LOANIO1_I16 ;
wire \hps_io|border|gpio_inst~LOANIO1_I17 ;
wire \hps_io|border|gpio_inst~LOANIO1_I18 ;
wire \hps_io|border|gpio_inst~LOANIO1_I19 ;
wire \hps_io|border|gpio_inst~LOANIO1_I20 ;
wire \hps_io|border|gpio_inst~LOANIO1_I21 ;
wire \hps_io|border|gpio_inst~LOANIO1_I22 ;
wire \hps_io|border|gpio_inst~LOANIO1_I23 ;
wire \hps_io|border|gpio_inst~LOANIO1_I24 ;
wire \hps_io|border|gpio_inst~LOANIO1_I25 ;
wire \hps_io|border|gpio_inst~LOANIO1_I26 ;
wire \hps_io|border|gpio_inst~LOANIO1_I27 ;
wire \hps_io|border|gpio_inst~LOANIO1_I28 ;
wire \hps_io|border|gpio_inst~LOANIO2_I0 ;
wire \hps_io|border|gpio_inst~LOANIO2_I1 ;
wire \hps_io|border|gpio_inst~LOANIO2_I2 ;
wire \hps_io|border|gpio_inst~LOANIO2_I3 ;
wire \hps_io|border|gpio_inst~LOANIO2_I4 ;
wire \hps_io|border|gpio_inst~LOANIO2_I5 ;
wire \hps_io|border|gpio_inst~LOANIO2_I6 ;
wire \hps_io|border|gpio_inst~LOANIO2_I7 ;
wire \hps_io|border|gpio_inst~LOANIO2_I8 ;


soc_system_soc_system_hps_0_fpga_interfaces fpga_interfaces(
	.loanio_gpio_loanio0_oe({\fpga_interfaces|loanio_gpio_loanio0_oe[28] ,\fpga_interfaces|loanio_gpio_loanio0_oe[27] ,\fpga_interfaces|loanio_gpio_loanio0_oe[26] ,\fpga_interfaces|loanio_gpio_loanio0_oe[25] ,\fpga_interfaces|loanio_gpio_loanio0_oe[24] ,
\fpga_interfaces|loanio_gpio_loanio0_oe[23] ,\fpga_interfaces|loanio_gpio_loanio0_oe[22] ,\fpga_interfaces|loanio_gpio_loanio0_oe[21] ,\fpga_interfaces|loanio_gpio_loanio0_oe[20] ,\fpga_interfaces|loanio_gpio_loanio0_oe[19] ,
\fpga_interfaces|loanio_gpio_loanio0_oe[18] ,\fpga_interfaces|loanio_gpio_loanio0_oe[17] ,\fpga_interfaces|loanio_gpio_loanio0_oe[16] ,\fpga_interfaces|loanio_gpio_loanio0_oe[15] ,\fpga_interfaces|loanio_gpio_loanio0_oe[14] ,
\fpga_interfaces|loanio_gpio_loanio0_oe[13] ,\fpga_interfaces|loanio_gpio_loanio0_oe[12] ,\fpga_interfaces|loanio_gpio_loanio0_oe[11] ,\fpga_interfaces|loanio_gpio_loanio0_oe[10] ,\fpga_interfaces|loanio_gpio_loanio0_oe[9] ,
\fpga_interfaces|loanio_gpio_loanio0_oe[8] ,\fpga_interfaces|loanio_gpio_loanio0_oe[7] ,\fpga_interfaces|loanio_gpio_loanio0_oe[6] ,\fpga_interfaces|loanio_gpio_loanio0_oe[5] ,\fpga_interfaces|loanio_gpio_loanio0_oe[4] ,
\fpga_interfaces|loanio_gpio_loanio0_oe[3] ,\fpga_interfaces|loanio_gpio_loanio0_oe[2] ,\fpga_interfaces|loanio_gpio_loanio0_oe[1] ,\fpga_interfaces|loanio_gpio_loanio0_oe[0] }),
	.loanio_gpio_loanio1_oe({\fpga_interfaces|loanio_gpio_loanio1_oe[28] ,\fpga_interfaces|loanio_gpio_loanio1_oe[27] ,\fpga_interfaces|loanio_gpio_loanio1_oe[26] ,\fpga_interfaces|loanio_gpio_loanio1_oe[25] ,\fpga_interfaces|loanio_gpio_loanio1_oe[24] ,
\fpga_interfaces|loanio_gpio_loanio1_oe[23] ,\fpga_interfaces|loanio_gpio_loanio1_oe[22] ,\fpga_interfaces|loanio_gpio_loanio1_oe[21] ,\fpga_interfaces|loanio_gpio_loanio1_oe[20] ,\fpga_interfaces|loanio_gpio_loanio1_oe[19] ,
\fpga_interfaces|loanio_gpio_loanio1_oe[18] ,\fpga_interfaces|loanio_gpio_loanio1_oe[17] ,\fpga_interfaces|loanio_gpio_loanio1_oe[16] ,\fpga_interfaces|loanio_gpio_loanio1_oe[15] ,\fpga_interfaces|loanio_gpio_loanio1_oe[14] ,
\fpga_interfaces|loanio_gpio_loanio1_oe[13] ,\fpga_interfaces|loanio_gpio_loanio1_oe[12] ,\fpga_interfaces|loanio_gpio_loanio1_oe[11] ,\fpga_interfaces|loanio_gpio_loanio1_oe[10] ,\fpga_interfaces|loanio_gpio_loanio1_oe[9] ,
\fpga_interfaces|loanio_gpio_loanio1_oe[8] ,\fpga_interfaces|loanio_gpio_loanio1_oe[7] ,\fpga_interfaces|loanio_gpio_loanio1_oe[6] ,\fpga_interfaces|loanio_gpio_loanio1_oe[5] ,\fpga_interfaces|loanio_gpio_loanio1_oe[4] ,
\fpga_interfaces|loanio_gpio_loanio1_oe[3] ,\fpga_interfaces|loanio_gpio_loanio1_oe[2] ,\fpga_interfaces|loanio_gpio_loanio1_oe[1] ,\fpga_interfaces|loanio_gpio_loanio1_oe[0] }),
	.loanio_gpio_loanio2_oe({\fpga_interfaces|loanio_gpio_loanio2_oe[8] ,\fpga_interfaces|loanio_gpio_loanio2_oe[7] ,\fpga_interfaces|loanio_gpio_loanio2_oe[6] ,\fpga_interfaces|loanio_gpio_loanio2_oe[5] ,\fpga_interfaces|loanio_gpio_loanio2_oe[4] ,
\fpga_interfaces|loanio_gpio_loanio2_oe[3] ,\fpga_interfaces|loanio_gpio_loanio2_oe[2] ,\fpga_interfaces|loanio_gpio_loanio2_oe[1] ,\fpga_interfaces|loanio_gpio_loanio2_oe[0] }),
	.loanio_gpio_loanio0_o({\fpga_interfaces|loanio_gpio_loanio0_o[28] ,\fpga_interfaces|loanio_gpio_loanio0_o[27] ,\fpga_interfaces|loanio_gpio_loanio0_o[26] ,\fpga_interfaces|loanio_gpio_loanio0_o[25] ,\fpga_interfaces|loanio_gpio_loanio0_o[24] ,
\fpga_interfaces|loanio_gpio_loanio0_o[23] ,\fpga_interfaces|loanio_gpio_loanio0_o[22] ,\fpga_interfaces|loanio_gpio_loanio0_o[21] ,\fpga_interfaces|loanio_gpio_loanio0_o[20] ,\fpga_interfaces|loanio_gpio_loanio0_o[19] ,
\fpga_interfaces|loanio_gpio_loanio0_o[18] ,\fpga_interfaces|loanio_gpio_loanio0_o[17] ,\fpga_interfaces|loanio_gpio_loanio0_o[16] ,\fpga_interfaces|loanio_gpio_loanio0_o[15] ,\fpga_interfaces|loanio_gpio_loanio0_o[14] ,
\fpga_interfaces|loanio_gpio_loanio0_o[13] ,\fpga_interfaces|loanio_gpio_loanio0_o[12] ,\fpga_interfaces|loanio_gpio_loanio0_o[11] ,\fpga_interfaces|loanio_gpio_loanio0_o[10] ,\fpga_interfaces|loanio_gpio_loanio0_o[9] ,\fpga_interfaces|loanio_gpio_loanio0_o[8] ,
\fpga_interfaces|loanio_gpio_loanio0_o[7] ,\fpga_interfaces|loanio_gpio_loanio0_o[6] ,\fpga_interfaces|loanio_gpio_loanio0_o[5] ,\fpga_interfaces|loanio_gpio_loanio0_o[4] ,\fpga_interfaces|loanio_gpio_loanio0_o[3] ,\fpga_interfaces|loanio_gpio_loanio0_o[2] ,
\fpga_interfaces|loanio_gpio_loanio0_o[1] ,\fpga_interfaces|loanio_gpio_loanio0_o[0] }),
	.loanio_gpio_loanio1_o({\fpga_interfaces|loanio_gpio_loanio1_o[28] ,\fpga_interfaces|loanio_gpio_loanio1_o[27] ,\fpga_interfaces|loanio_gpio_loanio1_o[26] ,\fpga_interfaces|loanio_gpio_loanio1_o[25] ,\fpga_interfaces|loanio_gpio_loanio1_o[24] ,
\fpga_interfaces|loanio_gpio_loanio1_o[23] ,\fpga_interfaces|loanio_gpio_loanio1_o[22] ,\fpga_interfaces|loanio_gpio_loanio1_o[21] ,\fpga_interfaces|loanio_gpio_loanio1_o[20] ,\fpga_interfaces|loanio_gpio_loanio1_o[19] ,
\fpga_interfaces|loanio_gpio_loanio1_o[18] ,\fpga_interfaces|loanio_gpio_loanio1_o[17] ,\fpga_interfaces|loanio_gpio_loanio1_o[16] ,\fpga_interfaces|loanio_gpio_loanio1_o[15] ,\fpga_interfaces|loanio_gpio_loanio1_o[14] ,
\fpga_interfaces|loanio_gpio_loanio1_o[13] ,\fpga_interfaces|loanio_gpio_loanio1_o[12] ,\fpga_interfaces|loanio_gpio_loanio1_o[11] ,\fpga_interfaces|loanio_gpio_loanio1_o[10] ,\fpga_interfaces|loanio_gpio_loanio1_o[9] ,\fpga_interfaces|loanio_gpio_loanio1_o[8] ,
\fpga_interfaces|loanio_gpio_loanio1_o[7] ,\fpga_interfaces|loanio_gpio_loanio1_o[6] ,\fpga_interfaces|loanio_gpio_loanio1_o[5] ,\fpga_interfaces|loanio_gpio_loanio1_o[4] ,\fpga_interfaces|loanio_gpio_loanio1_o[3] ,\fpga_interfaces|loanio_gpio_loanio1_o[2] ,
\fpga_interfaces|loanio_gpio_loanio1_o[1] ,\fpga_interfaces|loanio_gpio_loanio1_o[0] }),
	.loanio_gpio_loanio2_o({\fpga_interfaces|loanio_gpio_loanio2_o[8] ,\fpga_interfaces|loanio_gpio_loanio2_o[7] ,\fpga_interfaces|loanio_gpio_loanio2_o[6] ,\fpga_interfaces|loanio_gpio_loanio2_o[5] ,\fpga_interfaces|loanio_gpio_loanio2_o[4] ,\fpga_interfaces|loanio_gpio_loanio2_o[3] ,
\fpga_interfaces|loanio_gpio_loanio2_o[2] ,\fpga_interfaces|loanio_gpio_loanio2_o[1] ,\fpga_interfaces|loanio_gpio_loanio2_o[0] }),
	.h2f_loan_in({h2f_loan_in_66,h2f_loan_in_65,h2f_loan_in_64,h2f_loan_in_63,h2f_loan_in_62,h2f_loan_in_61,h2f_loan_in_60,h2f_loan_in_59,h2f_loan_in_58,h2f_loan_in_57,h2f_loan_in_56,h2f_loan_in_55,h2f_loan_in_54,h2f_loan_in_53,h2f_loan_in_52,h2f_loan_in_51,h2f_loan_in_50,h2f_loan_in_49,
h2f_loan_in_48,h2f_loan_in_47,h2f_loan_in_46,h2f_loan_in_45,h2f_loan_in_44,h2f_loan_in_43,h2f_loan_in_42,h2f_loan_in_41,h2f_loan_in_40,h2f_loan_in_39,h2f_loan_in_38,h2f_loan_in_37,h2f_loan_in_36,h2f_loan_in_35,h2f_loan_in_34,h2f_loan_in_33,h2f_loan_in_32,h2f_loan_in_31,
h2f_loan_in_30,h2f_loan_in_29,h2f_loan_in_28,h2f_loan_in_27,h2f_loan_in_26,h2f_loan_in_25,h2f_loan_in_24,h2f_loan_in_23,h2f_loan_in_22,h2f_loan_in_21,h2f_loan_in_20,h2f_loan_in_19,h2f_loan_in_18,h2f_loan_in_17,h2f_loan_in_16,h2f_loan_in_15,h2f_loan_in_14,h2f_loan_in_13,
h2f_loan_in_12,h2f_loan_in_11,h2f_loan_in_10,h2f_loan_in_9,h2f_loan_in_8,h2f_loan_in_7,h2f_loan_in_6,h2f_loan_in_5,h2f_loan_in_4,h2f_loan_in_3,h2f_loan_in_2,h2f_loan_in_1,h2f_loan_in_0}),
	.h2f_rst_n({h2f_rst_n_0}),
	.h2f_lw_ARVALID({h2f_lw_ARVALID_0}),
	.h2f_lw_AWVALID({h2f_lw_AWVALID_0}),
	.h2f_lw_BREADY({h2f_lw_BREADY_0}),
	.h2f_lw_RREADY({h2f_lw_RREADY_0}),
	.h2f_lw_WLAST({h2f_lw_WLAST_0}),
	.h2f_lw_WVALID({h2f_lw_WVALID_0}),
	.h2f_lw_ARADDR({h2f_lw_ARADDR_unconnected_wire_20,h2f_lw_ARADDR_unconnected_wire_19,h2f_lw_ARADDR_unconnected_wire_18,h2f_lw_ARADDR_unconnected_wire_17,h2f_lw_ARADDR_unconnected_wire_16,h2f_lw_ARADDR_unconnected_wire_15,h2f_lw_ARADDR_14,h2f_lw_ARADDR_13,h2f_lw_ARADDR_12,
h2f_lw_ARADDR_11,h2f_lw_ARADDR_10,h2f_lw_ARADDR_9,h2f_lw_ARADDR_8,h2f_lw_ARADDR_7,h2f_lw_ARADDR_6,h2f_lw_ARADDR_5,h2f_lw_ARADDR_4,h2f_lw_ARADDR_3,h2f_lw_ARADDR_2,h2f_lw_ARADDR_1,h2f_lw_ARADDR_0}),
	.h2f_lw_ARBURST({h2f_lw_ARBURST_1,h2f_lw_ARBURST_0}),
	.h2f_lw_ARID({h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0}),
	.h2f_lw_ARLEN({h2f_lw_ARLEN_3,h2f_lw_ARLEN_2,h2f_lw_ARLEN_1,h2f_lw_ARLEN_0}),
	.h2f_lw_ARSIZE({h2f_lw_ARSIZE_2,h2f_lw_ARSIZE_1,h2f_lw_ARSIZE_0}),
	.h2f_lw_AWADDR({h2f_lw_AWADDR_unconnected_wire_20,h2f_lw_AWADDR_unconnected_wire_19,h2f_lw_AWADDR_unconnected_wire_18,h2f_lw_AWADDR_unconnected_wire_17,h2f_lw_AWADDR_unconnected_wire_16,h2f_lw_AWADDR_unconnected_wire_15,h2f_lw_AWADDR_14,h2f_lw_AWADDR_13,h2f_lw_AWADDR_12,
h2f_lw_AWADDR_11,h2f_lw_AWADDR_10,h2f_lw_AWADDR_9,h2f_lw_AWADDR_8,h2f_lw_AWADDR_7,h2f_lw_AWADDR_6,h2f_lw_AWADDR_5,h2f_lw_AWADDR_4,h2f_lw_AWADDR_3,h2f_lw_AWADDR_2,h2f_lw_AWADDR_1,h2f_lw_AWADDR_0}),
	.h2f_lw_AWBURST({h2f_lw_AWBURST_1,h2f_lw_AWBURST_0}),
	.h2f_lw_AWID({h2f_lw_AWID_11,h2f_lw_AWID_10,h2f_lw_AWID_9,h2f_lw_AWID_8,h2f_lw_AWID_7,h2f_lw_AWID_6,h2f_lw_AWID_5,h2f_lw_AWID_4,h2f_lw_AWID_3,h2f_lw_AWID_2,h2f_lw_AWID_1,h2f_lw_AWID_0}),
	.h2f_lw_AWLEN({h2f_lw_AWLEN_3,h2f_lw_AWLEN_2,h2f_lw_AWLEN_1,h2f_lw_AWLEN_0}),
	.h2f_lw_AWSIZE({h2f_lw_AWSIZE_2,h2f_lw_AWSIZE_1,h2f_lw_AWSIZE_0}),
	.h2f_lw_WDATA({h2f_lw_WDATA_31,h2f_lw_WDATA_30,h2f_lw_WDATA_29,h2f_lw_WDATA_28,h2f_lw_WDATA_27,h2f_lw_WDATA_26,h2f_lw_WDATA_25,h2f_lw_WDATA_24,h2f_lw_WDATA_23,h2f_lw_WDATA_22,h2f_lw_WDATA_21,h2f_lw_WDATA_20,h2f_lw_WDATA_19,h2f_lw_WDATA_18,h2f_lw_WDATA_17,h2f_lw_WDATA_16,h2f_lw_WDATA_15,
h2f_lw_WDATA_14,h2f_lw_WDATA_13,h2f_lw_WDATA_12,h2f_lw_WDATA_11,h2f_lw_WDATA_10,h2f_lw_WDATA_9,h2f_lw_WDATA_8,h2f_lw_WDATA_7,h2f_lw_WDATA_6,h2f_lw_WDATA_5,h2f_lw_WDATA_4,h2f_lw_WDATA_3,h2f_lw_WDATA_2,h2f_lw_WDATA_1,h2f_lw_WDATA_0}),
	.h2f_lw_WSTRB({h2f_lw_WSTRB_3,h2f_lw_WSTRB_2,h2f_lw_WSTRB_1,h2f_lw_WSTRB_0}),
	.h2f_lw_axi_clk({outclk_wire_0}),
	.h2f_lw_ARREADY({sink1_ready}),
	.h2f_lw_AWREADY({awready}),
	.h2f_lw_BVALID({src0_valid}),
	.h2f_lw_RLAST({source_endofpacket}),
	.h2f_lw_RVALID({src1_valid}),
	.h2f_lw_WREADY({wready}),
	.h2f_lw_BID({mem_99_0,mem_98_0,mem_97_0,mem_96_0,mem_95_0,mem_94_0,mem_93_0,mem_92_0,mem_91_0,mem_90_0,mem_89_0,mem_88_0}),
	.h2f_lw_RID({mem_99_0,mem_98_0,mem_97_0,mem_96_0,mem_95_0,mem_94_0,mem_93_0,mem_92_0,mem_91_0,mem_90_0,mem_89_0,mem_88_0}),
	.h2f_lw_RDATA({out_data_31,out_data_30,out_data_29,out_data_28,out_data_27,out_data_26,out_data_25,out_data_24,out_data_23,out_data_22,out_data_21,out_data_20,out_data_19,out_data_18,out_data_17,out_data_16,out_data_15,out_data_14,out_data_13,out_data_12,out_data_11,out_data_10,out_data_9,
out_data_8,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.loanio_gpio_loanio0_i({\hps_io|border|gpio_inst~LOANIO0_I28 ,\hps_io|border|gpio_inst~LOANIO0_I27 ,\hps_io|border|gpio_inst~LOANIO0_I26 ,\hps_io|border|gpio_inst~LOANIO0_I25 ,\hps_io|border|gpio_inst~LOANIO0_I24 ,\hps_io|border|gpio_inst~LOANIO0_I23 ,
\hps_io|border|gpio_inst~LOANIO0_I22 ,\hps_io|border|gpio_inst~LOANIO0_I21 ,\hps_io|border|gpio_inst~LOANIO0_I20 ,\hps_io|border|gpio_inst~LOANIO0_I19 ,\hps_io|border|gpio_inst~LOANIO0_I18 ,\hps_io|border|gpio_inst~LOANIO0_I17 ,
\hps_io|border|gpio_inst~LOANIO0_I16 ,\hps_io|border|gpio_inst~LOANIO0_I15 ,\hps_io|border|gpio_inst~LOANIO0_I14 ,\hps_io|border|gpio_inst~LOANIO0_I13 ,\hps_io|border|gpio_inst~LOANIO0_I12 ,\hps_io|border|gpio_inst~LOANIO0_I11 ,
\hps_io|border|gpio_inst~LOANIO0_I10 ,\hps_io|border|gpio_inst~LOANIO0_I9 ,\hps_io|border|gpio_inst~LOANIO0_I8 ,\hps_io|border|gpio_inst~LOANIO0_I7 ,\hps_io|border|gpio_inst~LOANIO0_I6 ,\hps_io|border|gpio_inst~LOANIO0_I5 ,\hps_io|border|gpio_inst~LOANIO0_I4 ,
\hps_io|border|gpio_inst~LOANIO0_I3 ,\hps_io|border|gpio_inst~LOANIO0_I2 ,\hps_io|border|gpio_inst~LOANIO0_I1 ,\hps_io|border|gpio_inst~LOANIO0_I0 }),
	.loanio_gpio_loanio1_i({\hps_io|border|gpio_inst~LOANIO1_I28 ,\hps_io|border|gpio_inst~LOANIO1_I27 ,\hps_io|border|gpio_inst~LOANIO1_I26 ,\hps_io|border|gpio_inst~LOANIO1_I25 ,\hps_io|border|gpio_inst~LOANIO1_I24 ,\hps_io|border|gpio_inst~LOANIO1_I23 ,
\hps_io|border|gpio_inst~LOANIO1_I22 ,\hps_io|border|gpio_inst~LOANIO1_I21 ,\hps_io|border|gpio_inst~LOANIO1_I20 ,\hps_io|border|gpio_inst~LOANIO1_I19 ,\hps_io|border|gpio_inst~LOANIO1_I18 ,\hps_io|border|gpio_inst~LOANIO1_I17 ,
\hps_io|border|gpio_inst~LOANIO1_I16 ,\hps_io|border|gpio_inst~LOANIO1_I15 ,\hps_io|border|gpio_inst~LOANIO1_I14 ,\hps_io|border|gpio_inst~LOANIO1_I13 ,\hps_io|border|gpio_inst~LOANIO1_I12 ,\hps_io|border|gpio_inst~LOANIO1_I11 ,
\hps_io|border|gpio_inst~LOANIO1_I10 ,\hps_io|border|gpio_inst~LOANIO1_I9 ,\hps_io|border|gpio_inst~LOANIO1_I8 ,\hps_io|border|gpio_inst~LOANIO1_I7 ,\hps_io|border|gpio_inst~LOANIO1_I6 ,\hps_io|border|gpio_inst~LOANIO1_I5 ,\hps_io|border|gpio_inst~LOANIO1_I4 ,
\hps_io|border|gpio_inst~LOANIO1_I3 ,\hps_io|border|gpio_inst~LOANIO1_I2 ,\hps_io|border|gpio_inst~LOANIO1_I1 ,\hps_io|border|gpio_inst~LOANIO1_I0 }),
	.loanio_gpio_loanio2_i({\hps_io|border|gpio_inst~LOANIO2_I8 ,\hps_io|border|gpio_inst~LOANIO2_I7 ,\hps_io|border|gpio_inst~LOANIO2_I6 ,\hps_io|border|gpio_inst~LOANIO2_I5 ,\hps_io|border|gpio_inst~LOANIO2_I4 ,\hps_io|border|gpio_inst~LOANIO2_I3 ,\hps_io|border|gpio_inst~LOANIO2_I2 ,
\hps_io|border|gpio_inst~LOANIO2_I1 ,\hps_io|border|gpio_inst~LOANIO2_I0 }),
	.h2f_loan_oe({d_out_oe_66,d_out_oe_65,d_out_oe_64,d_out_oe_63,d_out_oe_62,d_out_oe_61,d_out_oe_60,d_out_oe_59,d_out_oe_58,d_out_oe_57,d_out_oe_56,d_out_oe_55,d_out_oe_54,d_out_oe_53,d_out_oe_52,d_out_oe_51,d_out_oe_50,d_out_oe_49,d_out_oe_48,d_out_oe_47,d_out_oe_46,d_out_oe_45,d_out_oe_44,
d_out_oe_43,d_out_oe_42,d_out_oe_41,d_out_oe_40,d_out_oe_39,d_out_oe_38,d_out_oe_37,d_out_oe_36,d_out_oe_35,d_out_oe_34,d_out_oe_33,d_out_oe_32,d_out_oe_31,d_out_oe_30,d_out_oe_29,d_out_oe_28,d_out_oe_27,d_out_oe_26,d_out_oe_25,d_out_oe_24,d_out_oe_23,d_out_oe_22,d_out_oe_21,
d_out_oe_20,d_out_oe_19,d_out_oe_18,d_out_oe_17,d_out_oe_16,d_out_oe_15,d_out_oe_14,d_out_oe_13,d_out_oe_12,d_out_oe_11,d_out_oe_10,d_out_oe_9,d_out_oe_8,d_out_oe_7,d_out_oe_6,d_out_oe_5,d_out_oe_4,d_out_oe_3,d_out_oe_2,d_out_oe_1,d_out_oe_0}),
	.h2f_loan_out({d_out_out_66,d_out_out_65,d_out_out_64,d_out_out_63,d_out_out_62,d_out_out_61,d_out_out_60,d_out_out_59,d_out_out_58,d_out_out_57,d_out_out_56,d_out_out_55,d_out_out_54,d_out_out_53,d_out_out_52,d_out_out_51,d_out_out_50,d_out_out_49,d_out_out_48,d_out_out_47,d_out_out_46,
d_out_out_45,d_out_out_44,d_out_out_43,d_out_out_42,d_out_out_41,d_out_out_40,d_out_out_39,d_out_out_38,d_out_out_37,d_out_out_36,d_out_out_35,d_out_out_34,d_out_out_33,d_out_out_32,d_out_out_31,d_out_out_30,d_out_out_29,d_out_out_28,d_out_out_27,d_out_out_26,d_out_out_25,
d_out_out_24,d_out_out_23,d_out_out_22,d_out_out_21,d_out_out_20,d_out_out_19,d_out_out_18,d_out_out_17,d_out_out_16,d_out_out_15,d_out_out_14,d_out_out_13,d_out_out_12,d_out_out_11,d_out_out_10,d_out_out_9,d_out_out_8,d_out_out_7,d_out_out_6,d_out_out_5,d_out_out_4,
d_out_out_3,d_out_out_2,d_out_out_1,d_out_out_0}));

soc_system_soc_system_hps_0_hps_io hps_io(
	.loanio_gpio_loanio0_oe_0(\fpga_interfaces|loanio_gpio_loanio0_oe[0] ),
	.loanio_gpio_loanio0_oe_1(\fpga_interfaces|loanio_gpio_loanio0_oe[1] ),
	.loanio_gpio_loanio0_oe_2(\fpga_interfaces|loanio_gpio_loanio0_oe[2] ),
	.loanio_gpio_loanio0_oe_3(\fpga_interfaces|loanio_gpio_loanio0_oe[3] ),
	.loanio_gpio_loanio0_oe_4(\fpga_interfaces|loanio_gpio_loanio0_oe[4] ),
	.loanio_gpio_loanio0_oe_5(\fpga_interfaces|loanio_gpio_loanio0_oe[5] ),
	.loanio_gpio_loanio0_oe_6(\fpga_interfaces|loanio_gpio_loanio0_oe[6] ),
	.loanio_gpio_loanio0_oe_7(\fpga_interfaces|loanio_gpio_loanio0_oe[7] ),
	.loanio_gpio_loanio0_oe_8(\fpga_interfaces|loanio_gpio_loanio0_oe[8] ),
	.loanio_gpio_loanio0_oe_9(\fpga_interfaces|loanio_gpio_loanio0_oe[9] ),
	.loanio_gpio_loanio0_oe_10(\fpga_interfaces|loanio_gpio_loanio0_oe[10] ),
	.loanio_gpio_loanio0_oe_11(\fpga_interfaces|loanio_gpio_loanio0_oe[11] ),
	.loanio_gpio_loanio0_oe_12(\fpga_interfaces|loanio_gpio_loanio0_oe[12] ),
	.loanio_gpio_loanio0_oe_13(\fpga_interfaces|loanio_gpio_loanio0_oe[13] ),
	.loanio_gpio_loanio0_oe_14(\fpga_interfaces|loanio_gpio_loanio0_oe[14] ),
	.loanio_gpio_loanio0_oe_15(\fpga_interfaces|loanio_gpio_loanio0_oe[15] ),
	.loanio_gpio_loanio0_oe_16(\fpga_interfaces|loanio_gpio_loanio0_oe[16] ),
	.loanio_gpio_loanio0_oe_17(\fpga_interfaces|loanio_gpio_loanio0_oe[17] ),
	.loanio_gpio_loanio0_oe_18(\fpga_interfaces|loanio_gpio_loanio0_oe[18] ),
	.loanio_gpio_loanio0_oe_19(\fpga_interfaces|loanio_gpio_loanio0_oe[19] ),
	.loanio_gpio_loanio0_oe_20(\fpga_interfaces|loanio_gpio_loanio0_oe[20] ),
	.loanio_gpio_loanio0_oe_21(\fpga_interfaces|loanio_gpio_loanio0_oe[21] ),
	.loanio_gpio_loanio0_oe_22(\fpga_interfaces|loanio_gpio_loanio0_oe[22] ),
	.loanio_gpio_loanio0_oe_23(\fpga_interfaces|loanio_gpio_loanio0_oe[23] ),
	.loanio_gpio_loanio0_oe_24(\fpga_interfaces|loanio_gpio_loanio0_oe[24] ),
	.loanio_gpio_loanio0_oe_25(\fpga_interfaces|loanio_gpio_loanio0_oe[25] ),
	.loanio_gpio_loanio0_oe_26(\fpga_interfaces|loanio_gpio_loanio0_oe[26] ),
	.loanio_gpio_loanio0_oe_27(\fpga_interfaces|loanio_gpio_loanio0_oe[27] ),
	.loanio_gpio_loanio0_oe_28(\fpga_interfaces|loanio_gpio_loanio0_oe[28] ),
	.loanio_gpio_loanio1_oe_0(\fpga_interfaces|loanio_gpio_loanio1_oe[0] ),
	.loanio_gpio_loanio1_oe_1(\fpga_interfaces|loanio_gpio_loanio1_oe[1] ),
	.loanio_gpio_loanio1_oe_2(\fpga_interfaces|loanio_gpio_loanio1_oe[2] ),
	.loanio_gpio_loanio1_oe_3(\fpga_interfaces|loanio_gpio_loanio1_oe[3] ),
	.loanio_gpio_loanio1_oe_4(\fpga_interfaces|loanio_gpio_loanio1_oe[4] ),
	.loanio_gpio_loanio1_oe_5(\fpga_interfaces|loanio_gpio_loanio1_oe[5] ),
	.loanio_gpio_loanio1_oe_6(\fpga_interfaces|loanio_gpio_loanio1_oe[6] ),
	.loanio_gpio_loanio1_oe_7(\fpga_interfaces|loanio_gpio_loanio1_oe[7] ),
	.loanio_gpio_loanio1_oe_8(\fpga_interfaces|loanio_gpio_loanio1_oe[8] ),
	.loanio_gpio_loanio1_oe_9(\fpga_interfaces|loanio_gpio_loanio1_oe[9] ),
	.loanio_gpio_loanio1_oe_10(\fpga_interfaces|loanio_gpio_loanio1_oe[10] ),
	.loanio_gpio_loanio1_oe_11(\fpga_interfaces|loanio_gpio_loanio1_oe[11] ),
	.loanio_gpio_loanio1_oe_12(\fpga_interfaces|loanio_gpio_loanio1_oe[12] ),
	.loanio_gpio_loanio1_oe_13(\fpga_interfaces|loanio_gpio_loanio1_oe[13] ),
	.loanio_gpio_loanio1_oe_14(\fpga_interfaces|loanio_gpio_loanio1_oe[14] ),
	.loanio_gpio_loanio1_oe_15(\fpga_interfaces|loanio_gpio_loanio1_oe[15] ),
	.loanio_gpio_loanio1_oe_16(\fpga_interfaces|loanio_gpio_loanio1_oe[16] ),
	.loanio_gpio_loanio1_oe_17(\fpga_interfaces|loanio_gpio_loanio1_oe[17] ),
	.loanio_gpio_loanio1_oe_18(\fpga_interfaces|loanio_gpio_loanio1_oe[18] ),
	.loanio_gpio_loanio1_oe_19(\fpga_interfaces|loanio_gpio_loanio1_oe[19] ),
	.loanio_gpio_loanio1_oe_20(\fpga_interfaces|loanio_gpio_loanio1_oe[20] ),
	.loanio_gpio_loanio1_oe_21(\fpga_interfaces|loanio_gpio_loanio1_oe[21] ),
	.loanio_gpio_loanio1_oe_22(\fpga_interfaces|loanio_gpio_loanio1_oe[22] ),
	.loanio_gpio_loanio1_oe_23(\fpga_interfaces|loanio_gpio_loanio1_oe[23] ),
	.loanio_gpio_loanio1_oe_24(\fpga_interfaces|loanio_gpio_loanio1_oe[24] ),
	.loanio_gpio_loanio1_oe_25(\fpga_interfaces|loanio_gpio_loanio1_oe[25] ),
	.loanio_gpio_loanio1_oe_26(\fpga_interfaces|loanio_gpio_loanio1_oe[26] ),
	.loanio_gpio_loanio1_oe_27(\fpga_interfaces|loanio_gpio_loanio1_oe[27] ),
	.loanio_gpio_loanio1_oe_28(\fpga_interfaces|loanio_gpio_loanio1_oe[28] ),
	.loanio_gpio_loanio2_oe_0(\fpga_interfaces|loanio_gpio_loanio2_oe[0] ),
	.loanio_gpio_loanio2_oe_1(\fpga_interfaces|loanio_gpio_loanio2_oe[1] ),
	.loanio_gpio_loanio2_oe_2(\fpga_interfaces|loanio_gpio_loanio2_oe[2] ),
	.loanio_gpio_loanio2_oe_3(\fpga_interfaces|loanio_gpio_loanio2_oe[3] ),
	.loanio_gpio_loanio2_oe_4(\fpga_interfaces|loanio_gpio_loanio2_oe[4] ),
	.loanio_gpio_loanio2_oe_5(\fpga_interfaces|loanio_gpio_loanio2_oe[5] ),
	.loanio_gpio_loanio2_oe_6(\fpga_interfaces|loanio_gpio_loanio2_oe[6] ),
	.loanio_gpio_loanio2_oe_7(\fpga_interfaces|loanio_gpio_loanio2_oe[7] ),
	.loanio_gpio_loanio2_oe_8(\fpga_interfaces|loanio_gpio_loanio2_oe[8] ),
	.loanio_gpio_loanio0_o_0(\fpga_interfaces|loanio_gpio_loanio0_o[0] ),
	.loanio_gpio_loanio0_o_1(\fpga_interfaces|loanio_gpio_loanio0_o[1] ),
	.loanio_gpio_loanio0_o_2(\fpga_interfaces|loanio_gpio_loanio0_o[2] ),
	.loanio_gpio_loanio0_o_3(\fpga_interfaces|loanio_gpio_loanio0_o[3] ),
	.loanio_gpio_loanio0_o_4(\fpga_interfaces|loanio_gpio_loanio0_o[4] ),
	.loanio_gpio_loanio0_o_5(\fpga_interfaces|loanio_gpio_loanio0_o[5] ),
	.loanio_gpio_loanio0_o_6(\fpga_interfaces|loanio_gpio_loanio0_o[6] ),
	.loanio_gpio_loanio0_o_7(\fpga_interfaces|loanio_gpio_loanio0_o[7] ),
	.loanio_gpio_loanio0_o_8(\fpga_interfaces|loanio_gpio_loanio0_o[8] ),
	.loanio_gpio_loanio0_o_9(\fpga_interfaces|loanio_gpio_loanio0_o[9] ),
	.loanio_gpio_loanio0_o_10(\fpga_interfaces|loanio_gpio_loanio0_o[10] ),
	.loanio_gpio_loanio0_o_11(\fpga_interfaces|loanio_gpio_loanio0_o[11] ),
	.loanio_gpio_loanio0_o_12(\fpga_interfaces|loanio_gpio_loanio0_o[12] ),
	.loanio_gpio_loanio0_o_13(\fpga_interfaces|loanio_gpio_loanio0_o[13] ),
	.loanio_gpio_loanio0_o_14(\fpga_interfaces|loanio_gpio_loanio0_o[14] ),
	.loanio_gpio_loanio0_o_15(\fpga_interfaces|loanio_gpio_loanio0_o[15] ),
	.loanio_gpio_loanio0_o_16(\fpga_interfaces|loanio_gpio_loanio0_o[16] ),
	.loanio_gpio_loanio0_o_17(\fpga_interfaces|loanio_gpio_loanio0_o[17] ),
	.loanio_gpio_loanio0_o_18(\fpga_interfaces|loanio_gpio_loanio0_o[18] ),
	.loanio_gpio_loanio0_o_19(\fpga_interfaces|loanio_gpio_loanio0_o[19] ),
	.loanio_gpio_loanio0_o_20(\fpga_interfaces|loanio_gpio_loanio0_o[20] ),
	.loanio_gpio_loanio0_o_21(\fpga_interfaces|loanio_gpio_loanio0_o[21] ),
	.loanio_gpio_loanio0_o_22(\fpga_interfaces|loanio_gpio_loanio0_o[22] ),
	.loanio_gpio_loanio0_o_23(\fpga_interfaces|loanio_gpio_loanio0_o[23] ),
	.loanio_gpio_loanio0_o_24(\fpga_interfaces|loanio_gpio_loanio0_o[24] ),
	.loanio_gpio_loanio0_o_25(\fpga_interfaces|loanio_gpio_loanio0_o[25] ),
	.loanio_gpio_loanio0_o_26(\fpga_interfaces|loanio_gpio_loanio0_o[26] ),
	.loanio_gpio_loanio0_o_27(\fpga_interfaces|loanio_gpio_loanio0_o[27] ),
	.loanio_gpio_loanio0_o_28(\fpga_interfaces|loanio_gpio_loanio0_o[28] ),
	.loanio_gpio_loanio1_o_0(\fpga_interfaces|loanio_gpio_loanio1_o[0] ),
	.loanio_gpio_loanio1_o_1(\fpga_interfaces|loanio_gpio_loanio1_o[1] ),
	.loanio_gpio_loanio1_o_2(\fpga_interfaces|loanio_gpio_loanio1_o[2] ),
	.loanio_gpio_loanio1_o_3(\fpga_interfaces|loanio_gpio_loanio1_o[3] ),
	.loanio_gpio_loanio1_o_4(\fpga_interfaces|loanio_gpio_loanio1_o[4] ),
	.loanio_gpio_loanio1_o_5(\fpga_interfaces|loanio_gpio_loanio1_o[5] ),
	.loanio_gpio_loanio1_o_6(\fpga_interfaces|loanio_gpio_loanio1_o[6] ),
	.loanio_gpio_loanio1_o_7(\fpga_interfaces|loanio_gpio_loanio1_o[7] ),
	.loanio_gpio_loanio1_o_8(\fpga_interfaces|loanio_gpio_loanio1_o[8] ),
	.loanio_gpio_loanio1_o_9(\fpga_interfaces|loanio_gpio_loanio1_o[9] ),
	.loanio_gpio_loanio1_o_10(\fpga_interfaces|loanio_gpio_loanio1_o[10] ),
	.loanio_gpio_loanio1_o_11(\fpga_interfaces|loanio_gpio_loanio1_o[11] ),
	.loanio_gpio_loanio1_o_12(\fpga_interfaces|loanio_gpio_loanio1_o[12] ),
	.loanio_gpio_loanio1_o_13(\fpga_interfaces|loanio_gpio_loanio1_o[13] ),
	.loanio_gpio_loanio1_o_14(\fpga_interfaces|loanio_gpio_loanio1_o[14] ),
	.loanio_gpio_loanio1_o_15(\fpga_interfaces|loanio_gpio_loanio1_o[15] ),
	.loanio_gpio_loanio1_o_16(\fpga_interfaces|loanio_gpio_loanio1_o[16] ),
	.loanio_gpio_loanio1_o_17(\fpga_interfaces|loanio_gpio_loanio1_o[17] ),
	.loanio_gpio_loanio1_o_18(\fpga_interfaces|loanio_gpio_loanio1_o[18] ),
	.loanio_gpio_loanio1_o_19(\fpga_interfaces|loanio_gpio_loanio1_o[19] ),
	.loanio_gpio_loanio1_o_20(\fpga_interfaces|loanio_gpio_loanio1_o[20] ),
	.loanio_gpio_loanio1_o_21(\fpga_interfaces|loanio_gpio_loanio1_o[21] ),
	.loanio_gpio_loanio1_o_22(\fpga_interfaces|loanio_gpio_loanio1_o[22] ),
	.loanio_gpio_loanio1_o_23(\fpga_interfaces|loanio_gpio_loanio1_o[23] ),
	.loanio_gpio_loanio1_o_24(\fpga_interfaces|loanio_gpio_loanio1_o[24] ),
	.loanio_gpio_loanio1_o_25(\fpga_interfaces|loanio_gpio_loanio1_o[25] ),
	.loanio_gpio_loanio1_o_26(\fpga_interfaces|loanio_gpio_loanio1_o[26] ),
	.loanio_gpio_loanio1_o_27(\fpga_interfaces|loanio_gpio_loanio1_o[27] ),
	.loanio_gpio_loanio1_o_28(\fpga_interfaces|loanio_gpio_loanio1_o[28] ),
	.loanio_gpio_loanio2_o_0(\fpga_interfaces|loanio_gpio_loanio2_o[0] ),
	.loanio_gpio_loanio2_o_1(\fpga_interfaces|loanio_gpio_loanio2_o[1] ),
	.loanio_gpio_loanio2_o_2(\fpga_interfaces|loanio_gpio_loanio2_o[2] ),
	.loanio_gpio_loanio2_o_3(\fpga_interfaces|loanio_gpio_loanio2_o[3] ),
	.loanio_gpio_loanio2_o_4(\fpga_interfaces|loanio_gpio_loanio2_o[4] ),
	.loanio_gpio_loanio2_o_5(\fpga_interfaces|loanio_gpio_loanio2_o[5] ),
	.loanio_gpio_loanio2_o_6(\fpga_interfaces|loanio_gpio_loanio2_o[6] ),
	.loanio_gpio_loanio2_o_7(\fpga_interfaces|loanio_gpio_loanio2_o[7] ),
	.loanio_gpio_loanio2_o_8(\fpga_interfaces|loanio_gpio_loanio2_o[8] ),
	.emac1_inst(emac1_inst),
	.emac1_inst1(emac1_inst1),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.emac1_inst2(emac1_inst2),
	.emac1_inst3(emac1_inst3),
	.emac1_inst4(emac1_inst4),
	.emac1_inst5(emac1_inst5),
	.emac1_inst6(emac1_inst6),
	.qspi_inst(qspi_inst),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.qspi_inst1(qspi_inst1),
	.sdio_inst(sdio_inst),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.usb1_inst(usb1_inst),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.spim0_inst(spim0_inst),
	.spim0_inst1(spim0_inst1),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.spim1_inst(spim1_inst),
	.spim1_inst1(spim1_inst1),
	.intermediate_38(intermediate_38),
	.intermediate_39(intermediate_39),
	.uart0_inst(uart0_inst),
	.gpio_inst(\hps_io|border|gpio_inst~LOANIO0_I0 ),
	.gpio_inst1(\hps_io|border|gpio_inst~LOANIO0_I1 ),
	.gpio_inst2(\hps_io|border|gpio_inst~LOANIO0_I2 ),
	.gpio_inst3(\hps_io|border|gpio_inst~LOANIO0_I3 ),
	.gpio_inst4(\hps_io|border|gpio_inst~LOANIO0_I4 ),
	.gpio_inst5(\hps_io|border|gpio_inst~LOANIO0_I5 ),
	.gpio_inst6(\hps_io|border|gpio_inst~LOANIO0_I6 ),
	.gpio_inst7(\hps_io|border|gpio_inst~LOANIO0_I7 ),
	.gpio_inst8(\hps_io|border|gpio_inst~LOANIO0_I8 ),
	.gpio_inst9(\hps_io|border|gpio_inst~LOANIO0_I9 ),
	.gpio_inst10(\hps_io|border|gpio_inst~LOANIO0_I10 ),
	.gpio_inst11(\hps_io|border|gpio_inst~LOANIO0_I11 ),
	.gpio_inst12(\hps_io|border|gpio_inst~LOANIO0_I12 ),
	.gpio_inst13(\hps_io|border|gpio_inst~LOANIO0_I13 ),
	.gpio_inst14(\hps_io|border|gpio_inst~LOANIO0_I14 ),
	.gpio_inst15(\hps_io|border|gpio_inst~LOANIO0_I15 ),
	.gpio_inst16(\hps_io|border|gpio_inst~LOANIO0_I16 ),
	.gpio_inst17(\hps_io|border|gpio_inst~LOANIO0_I17 ),
	.gpio_inst18(\hps_io|border|gpio_inst~LOANIO0_I18 ),
	.gpio_inst19(\hps_io|border|gpio_inst~LOANIO0_I19 ),
	.gpio_inst20(\hps_io|border|gpio_inst~LOANIO0_I20 ),
	.gpio_inst21(\hps_io|border|gpio_inst~LOANIO0_I21 ),
	.gpio_inst22(\hps_io|border|gpio_inst~LOANIO0_I22 ),
	.gpio_inst23(\hps_io|border|gpio_inst~LOANIO0_I23 ),
	.gpio_inst24(\hps_io|border|gpio_inst~LOANIO0_I24 ),
	.gpio_inst25(\hps_io|border|gpio_inst~LOANIO0_I25 ),
	.gpio_inst26(\hps_io|border|gpio_inst~LOANIO0_I26 ),
	.gpio_inst27(\hps_io|border|gpio_inst~LOANIO0_I27 ),
	.gpio_inst28(\hps_io|border|gpio_inst~LOANIO0_I28 ),
	.gpio_inst29(\hps_io|border|gpio_inst~LOANIO1_I0 ),
	.gpio_inst30(\hps_io|border|gpio_inst~LOANIO1_I1 ),
	.gpio_inst31(\hps_io|border|gpio_inst~LOANIO1_I2 ),
	.gpio_inst32(\hps_io|border|gpio_inst~LOANIO1_I3 ),
	.gpio_inst33(\hps_io|border|gpio_inst~LOANIO1_I4 ),
	.gpio_inst34(\hps_io|border|gpio_inst~LOANIO1_I5 ),
	.gpio_inst35(\hps_io|border|gpio_inst~LOANIO1_I6 ),
	.gpio_inst36(\hps_io|border|gpio_inst~LOANIO1_I7 ),
	.gpio_inst37(\hps_io|border|gpio_inst~LOANIO1_I8 ),
	.gpio_inst38(\hps_io|border|gpio_inst~LOANIO1_I9 ),
	.gpio_inst39(\hps_io|border|gpio_inst~LOANIO1_I10 ),
	.gpio_inst40(\hps_io|border|gpio_inst~LOANIO1_I11 ),
	.gpio_inst41(\hps_io|border|gpio_inst~LOANIO1_I12 ),
	.gpio_inst42(\hps_io|border|gpio_inst~LOANIO1_I13 ),
	.gpio_inst43(\hps_io|border|gpio_inst~LOANIO1_I14 ),
	.gpio_inst44(\hps_io|border|gpio_inst~LOANIO1_I15 ),
	.gpio_inst45(\hps_io|border|gpio_inst~LOANIO1_I16 ),
	.gpio_inst46(\hps_io|border|gpio_inst~LOANIO1_I17 ),
	.gpio_inst47(\hps_io|border|gpio_inst~LOANIO1_I18 ),
	.gpio_inst48(\hps_io|border|gpio_inst~LOANIO1_I19 ),
	.gpio_inst49(\hps_io|border|gpio_inst~LOANIO1_I20 ),
	.gpio_inst50(\hps_io|border|gpio_inst~LOANIO1_I21 ),
	.gpio_inst51(\hps_io|border|gpio_inst~LOANIO1_I22 ),
	.gpio_inst52(\hps_io|border|gpio_inst~LOANIO1_I23 ),
	.gpio_inst53(\hps_io|border|gpio_inst~LOANIO1_I24 ),
	.gpio_inst54(\hps_io|border|gpio_inst~LOANIO1_I25 ),
	.gpio_inst55(\hps_io|border|gpio_inst~LOANIO1_I26 ),
	.gpio_inst56(\hps_io|border|gpio_inst~LOANIO1_I27 ),
	.gpio_inst57(\hps_io|border|gpio_inst~LOANIO1_I28 ),
	.gpio_inst58(\hps_io|border|gpio_inst~LOANIO2_I0 ),
	.gpio_inst59(\hps_io|border|gpio_inst~LOANIO2_I1 ),
	.gpio_inst60(\hps_io|border|gpio_inst~LOANIO2_I2 ),
	.gpio_inst61(\hps_io|border|gpio_inst~LOANIO2_I3 ),
	.gpio_inst62(\hps_io|border|gpio_inst~LOANIO2_I4 ),
	.gpio_inst63(\hps_io|border|gpio_inst~LOANIO2_I5 ),
	.gpio_inst64(\hps_io|border|gpio_inst~LOANIO2_I6 ),
	.gpio_inst65(\hps_io|border|gpio_inst~LOANIO2_I7 ),
	.gpio_inst66(\hps_io|border|gpio_inst~LOANIO2_I8 ),
	.intermediate_50(intermediate_50),
	.intermediate_40(intermediate_40),
	.intermediate_51(intermediate_51),
	.intermediate_41(intermediate_41),
	.intermediate_42(intermediate_42),
	.intermediate_52(intermediate_52),
	.intermediate_44(intermediate_44),
	.intermediate_54(intermediate_54),
	.intermediate_56(intermediate_56),
	.intermediate_58(intermediate_58),
	.intermediate_60(intermediate_60),
	.intermediate_62(intermediate_62),
	.intermediate_64(intermediate_64),
	.intermediate_43(intermediate_43),
	.intermediate_53(intermediate_53),
	.intermediate_45(intermediate_45),
	.intermediate_55(intermediate_55),
	.intermediate_57(intermediate_57),
	.intermediate_59(intermediate_59),
	.intermediate_61(intermediate_61),
	.intermediate_63(intermediate_63),
	.intermediate_65(intermediate_65),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_gpio_inst_GPIO62_0(hps_io_gpio_inst_GPIO62_0),
	.hps_io_gpio_inst_LOANIO00_0(hps_io_gpio_inst_LOANIO00_0),
	.hps_io_gpio_inst_LOANIO41_0(hps_io_gpio_inst_LOANIO41_0),
	.hps_io_gpio_inst_LOANIO51_0(hps_io_gpio_inst_LOANIO51_0),
	.hps_io_gpio_inst_LOANIO52_0(hps_io_gpio_inst_LOANIO52_0),
	.hps_io_gpio_inst_LOANIO53_0(hps_io_gpio_inst_LOANIO53_0),
	.hps_io_gpio_inst_LOANIO54_0(hps_io_gpio_inst_LOANIO54_0),
	.hps_io_gpio_inst_LOANIO55_0(hps_io_gpio_inst_LOANIO55_0),
	.hps_io_gpio_inst_LOANIO56_0(hps_io_gpio_inst_LOANIO56_0),
	.hps_io_hps_io_emac1_inst_RXD0(hps_io_hps_io_emac1_inst_RXD0),
	.hps_io_hps_io_emac1_inst_RXD1(hps_io_hps_io_emac1_inst_RXD1),
	.hps_io_hps_io_emac1_inst_RXD2(hps_io_hps_io_emac1_inst_RXD2),
	.hps_io_hps_io_emac1_inst_RXD3(hps_io_hps_io_emac1_inst_RXD3),
	.hps_io_hps_io_emac1_inst_RX_CLK(hps_io_hps_io_emac1_inst_RX_CLK),
	.hps_io_hps_io_emac1_inst_RX_CTL(hps_io_hps_io_emac1_inst_RX_CTL),
	.hps_io_hps_io_spim0_inst_MISO(hps_io_hps_io_spim0_inst_MISO),
	.hps_io_hps_io_spim1_inst_MISO(hps_io_hps_io_spim1_inst_MISO),
	.hps_io_hps_io_uart0_inst_RX(hps_io_hps_io_uart0_inst_RX),
	.hps_io_hps_io_usb1_inst_CLK(hps_io_hps_io_usb1_inst_CLK),
	.hps_io_hps_io_usb1_inst_DIR(hps_io_hps_io_usb1_inst_DIR),
	.hps_io_hps_io_usb1_inst_NXT(hps_io_hps_io_usb1_inst_NXT),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module soc_system_soc_system_hps_0_fpga_interfaces (
	loanio_gpio_loanio0_oe,
	loanio_gpio_loanio1_oe,
	loanio_gpio_loanio2_oe,
	loanio_gpio_loanio0_o,
	loanio_gpio_loanio1_o,
	loanio_gpio_loanio2_o,
	h2f_loan_in,
	h2f_rst_n,
	h2f_lw_ARVALID,
	h2f_lw_AWVALID,
	h2f_lw_BREADY,
	h2f_lw_RREADY,
	h2f_lw_WLAST,
	h2f_lw_WVALID,
	h2f_lw_ARADDR,
	h2f_lw_ARBURST,
	h2f_lw_ARID,
	h2f_lw_ARLEN,
	h2f_lw_ARSIZE,
	h2f_lw_AWADDR,
	h2f_lw_AWBURST,
	h2f_lw_AWID,
	h2f_lw_AWLEN,
	h2f_lw_AWSIZE,
	h2f_lw_WDATA,
	h2f_lw_WSTRB,
	h2f_lw_axi_clk,
	h2f_lw_ARREADY,
	h2f_lw_AWREADY,
	h2f_lw_BVALID,
	h2f_lw_RLAST,
	h2f_lw_RVALID,
	h2f_lw_WREADY,
	h2f_lw_BID,
	h2f_lw_RID,
	h2f_lw_RDATA,
	loanio_gpio_loanio0_i,
	loanio_gpio_loanio1_i,
	loanio_gpio_loanio2_i,
	h2f_loan_oe,
	h2f_loan_out)/* synthesis synthesis_greybox=0 */;
output 	[28:0] loanio_gpio_loanio0_oe;
output 	[28:0] loanio_gpio_loanio1_oe;
output 	[8:0] loanio_gpio_loanio2_oe;
output 	[28:0] loanio_gpio_loanio0_o;
output 	[28:0] loanio_gpio_loanio1_o;
output 	[8:0] loanio_gpio_loanio2_o;
output 	[66:0] h2f_loan_in;
output 	[0:0] h2f_rst_n;
output 	[0:0] h2f_lw_ARVALID;
output 	[0:0] h2f_lw_AWVALID;
output 	[0:0] h2f_lw_BREADY;
output 	[0:0] h2f_lw_RREADY;
output 	[0:0] h2f_lw_WLAST;
output 	[0:0] h2f_lw_WVALID;
output 	[20:0] h2f_lw_ARADDR;
output 	[1:0] h2f_lw_ARBURST;
output 	[11:0] h2f_lw_ARID;
output 	[3:0] h2f_lw_ARLEN;
output 	[2:0] h2f_lw_ARSIZE;
output 	[20:0] h2f_lw_AWADDR;
output 	[1:0] h2f_lw_AWBURST;
output 	[11:0] h2f_lw_AWID;
output 	[3:0] h2f_lw_AWLEN;
output 	[2:0] h2f_lw_AWSIZE;
output 	[31:0] h2f_lw_WDATA;
output 	[3:0] h2f_lw_WSTRB;
input 	[0:0] h2f_lw_axi_clk;
input 	[0:0] h2f_lw_ARREADY;
input 	[0:0] h2f_lw_AWREADY;
input 	[0:0] h2f_lw_BVALID;
input 	[0:0] h2f_lw_RLAST;
input 	[0:0] h2f_lw_RVALID;
input 	[0:0] h2f_lw_WREADY;
input 	[11:0] h2f_lw_BID;
input 	[11:0] h2f_lw_RID;
input 	[31:0] h2f_lw_RDATA;
input 	[28:0] loanio_gpio_loanio0_i;
input 	[28:0] loanio_gpio_loanio1_i;
input 	[8:0] loanio_gpio_loanio2_i;
input 	[66:0] h2f_loan_oe;
input 	[66:0] h2f_loan_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \fpga2hps~arready ;
wire \hps2fpga~araddr ;
wire \hps2fpga~O_ARADDR1 ;
wire \hps2fpga~O_ARADDR2 ;
wire \hps2fpga~O_ARADDR3 ;
wire \hps2fpga~O_ARADDR4 ;
wire \hps2fpga~O_ARADDR5 ;
wire \hps2fpga~O_ARADDR6 ;
wire \hps2fpga~O_ARADDR7 ;
wire \hps2fpga~O_ARADDR8 ;
wire \hps2fpga~O_ARADDR9 ;
wire \hps2fpga~O_ARADDR10 ;
wire \hps2fpga~O_ARADDR11 ;
wire \hps2fpga~O_ARADDR12 ;
wire \hps2fpga~O_ARADDR13 ;
wire \hps2fpga~O_ARADDR14 ;
wire \hps2fpga~O_ARADDR15 ;
wire \hps2fpga~O_ARADDR16 ;
wire \hps2fpga~O_ARADDR17 ;
wire \hps2fpga~O_ARADDR18 ;
wire \hps2fpga~O_ARADDR19 ;
wire \hps2fpga~O_ARADDR20 ;
wire \hps2fpga~O_ARADDR21 ;
wire \hps2fpga~O_ARADDR22 ;
wire \hps2fpga~O_ARADDR23 ;
wire \hps2fpga~O_ARADDR24 ;
wire \hps2fpga~O_ARADDR25 ;
wire \hps2fpga~O_ARADDR26 ;
wire \hps2fpga~O_ARADDR27 ;
wire \hps2fpga~O_ARADDR28 ;
wire \hps2fpga~O_ARADDR29 ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \loan_io_inst~fake_dout ;
wire \clocks_resets~h2f_cold_rst_n ;
wire \h2f_lw_ARADDR[15] ;
wire \h2f_lw_ARADDR[16] ;
wire \h2f_lw_ARADDR[17] ;
wire \h2f_lw_ARADDR[18] ;
wire \h2f_lw_ARADDR[19] ;
wire \h2f_lw_ARADDR[20] ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [70:0] loan_io_inst_GPIO_OE_bus;
wire [70:0] loan_io_inst_GPIO_OUT_bus;
wire [70:0] loan_io_inst_LOANIO_IN_bus;
wire [20:0] hps2fpga_light_weight_ARADDR_bus;
wire [1:0] hps2fpga_light_weight_ARBURST_bus;
wire [11:0] hps2fpga_light_weight_ARID_bus;
wire [3:0] hps2fpga_light_weight_ARLEN_bus;
wire [2:0] hps2fpga_light_weight_ARSIZE_bus;
wire [20:0] hps2fpga_light_weight_AWADDR_bus;
wire [1:0] hps2fpga_light_weight_AWBURST_bus;
wire [11:0] hps2fpga_light_weight_AWID_bus;
wire [3:0] hps2fpga_light_weight_AWLEN_bus;
wire [2:0] hps2fpga_light_weight_AWSIZE_bus;
wire [31:0] hps2fpga_light_weight_WDATA_bus;
wire [3:0] hps2fpga_light_weight_WSTRB_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \hps2fpga~araddr  = hps2fpga_ARADDR_bus[0];
assign \hps2fpga~O_ARADDR1  = hps2fpga_ARADDR_bus[1];
assign \hps2fpga~O_ARADDR2  = hps2fpga_ARADDR_bus[2];
assign \hps2fpga~O_ARADDR3  = hps2fpga_ARADDR_bus[3];
assign \hps2fpga~O_ARADDR4  = hps2fpga_ARADDR_bus[4];
assign \hps2fpga~O_ARADDR5  = hps2fpga_ARADDR_bus[5];
assign \hps2fpga~O_ARADDR6  = hps2fpga_ARADDR_bus[6];
assign \hps2fpga~O_ARADDR7  = hps2fpga_ARADDR_bus[7];
assign \hps2fpga~O_ARADDR8  = hps2fpga_ARADDR_bus[8];
assign \hps2fpga~O_ARADDR9  = hps2fpga_ARADDR_bus[9];
assign \hps2fpga~O_ARADDR10  = hps2fpga_ARADDR_bus[10];
assign \hps2fpga~O_ARADDR11  = hps2fpga_ARADDR_bus[11];
assign \hps2fpga~O_ARADDR12  = hps2fpga_ARADDR_bus[12];
assign \hps2fpga~O_ARADDR13  = hps2fpga_ARADDR_bus[13];
assign \hps2fpga~O_ARADDR14  = hps2fpga_ARADDR_bus[14];
assign \hps2fpga~O_ARADDR15  = hps2fpga_ARADDR_bus[15];
assign \hps2fpga~O_ARADDR16  = hps2fpga_ARADDR_bus[16];
assign \hps2fpga~O_ARADDR17  = hps2fpga_ARADDR_bus[17];
assign \hps2fpga~O_ARADDR18  = hps2fpga_ARADDR_bus[18];
assign \hps2fpga~O_ARADDR19  = hps2fpga_ARADDR_bus[19];
assign \hps2fpga~O_ARADDR20  = hps2fpga_ARADDR_bus[20];
assign \hps2fpga~O_ARADDR21  = hps2fpga_ARADDR_bus[21];
assign \hps2fpga~O_ARADDR22  = hps2fpga_ARADDR_bus[22];
assign \hps2fpga~O_ARADDR23  = hps2fpga_ARADDR_bus[23];
assign \hps2fpga~O_ARADDR24  = hps2fpga_ARADDR_bus[24];
assign \hps2fpga~O_ARADDR25  = hps2fpga_ARADDR_bus[25];
assign \hps2fpga~O_ARADDR26  = hps2fpga_ARADDR_bus[26];
assign \hps2fpga~O_ARADDR27  = hps2fpga_ARADDR_bus[27];
assign \hps2fpga~O_ARADDR28  = hps2fpga_ARADDR_bus[28];
assign \hps2fpga~O_ARADDR29  = hps2fpga_ARADDR_bus[29];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign loanio_gpio_loanio0_oe[0] = loan_io_inst_GPIO_OE_bus[0];
assign loanio_gpio_loanio0_oe[1] = loan_io_inst_GPIO_OE_bus[1];
assign loanio_gpio_loanio0_oe[2] = loan_io_inst_GPIO_OE_bus[2];
assign loanio_gpio_loanio0_oe[3] = loan_io_inst_GPIO_OE_bus[3];
assign loanio_gpio_loanio0_oe[4] = loan_io_inst_GPIO_OE_bus[4];
assign loanio_gpio_loanio0_oe[5] = loan_io_inst_GPIO_OE_bus[5];
assign loanio_gpio_loanio0_oe[6] = loan_io_inst_GPIO_OE_bus[6];
assign loanio_gpio_loanio0_oe[7] = loan_io_inst_GPIO_OE_bus[7];
assign loanio_gpio_loanio0_oe[8] = loan_io_inst_GPIO_OE_bus[8];
assign loanio_gpio_loanio0_oe[9] = loan_io_inst_GPIO_OE_bus[9];
assign loanio_gpio_loanio0_oe[10] = loan_io_inst_GPIO_OE_bus[10];
assign loanio_gpio_loanio0_oe[11] = loan_io_inst_GPIO_OE_bus[11];
assign loanio_gpio_loanio0_oe[12] = loan_io_inst_GPIO_OE_bus[12];
assign loanio_gpio_loanio0_oe[13] = loan_io_inst_GPIO_OE_bus[13];
assign loanio_gpio_loanio0_oe[14] = loan_io_inst_GPIO_OE_bus[14];
assign loanio_gpio_loanio0_oe[15] = loan_io_inst_GPIO_OE_bus[15];
assign loanio_gpio_loanio0_oe[16] = loan_io_inst_GPIO_OE_bus[16];
assign loanio_gpio_loanio0_oe[17] = loan_io_inst_GPIO_OE_bus[17];
assign loanio_gpio_loanio0_oe[18] = loan_io_inst_GPIO_OE_bus[18];
assign loanio_gpio_loanio0_oe[19] = loan_io_inst_GPIO_OE_bus[19];
assign loanio_gpio_loanio0_oe[20] = loan_io_inst_GPIO_OE_bus[20];
assign loanio_gpio_loanio0_oe[21] = loan_io_inst_GPIO_OE_bus[21];
assign loanio_gpio_loanio0_oe[22] = loan_io_inst_GPIO_OE_bus[22];
assign loanio_gpio_loanio0_oe[23] = loan_io_inst_GPIO_OE_bus[23];
assign loanio_gpio_loanio0_oe[24] = loan_io_inst_GPIO_OE_bus[24];
assign loanio_gpio_loanio0_oe[25] = loan_io_inst_GPIO_OE_bus[25];
assign loanio_gpio_loanio0_oe[26] = loan_io_inst_GPIO_OE_bus[26];
assign loanio_gpio_loanio0_oe[27] = loan_io_inst_GPIO_OE_bus[27];
assign loanio_gpio_loanio0_oe[28] = loan_io_inst_GPIO_OE_bus[28];
assign loanio_gpio_loanio1_oe[0] = loan_io_inst_GPIO_OE_bus[29];
assign loanio_gpio_loanio1_oe[1] = loan_io_inst_GPIO_OE_bus[30];
assign loanio_gpio_loanio1_oe[2] = loan_io_inst_GPIO_OE_bus[31];
assign loanio_gpio_loanio1_oe[3] = loan_io_inst_GPIO_OE_bus[32];
assign loanio_gpio_loanio1_oe[4] = loan_io_inst_GPIO_OE_bus[33];
assign loanio_gpio_loanio1_oe[5] = loan_io_inst_GPIO_OE_bus[34];
assign loanio_gpio_loanio1_oe[6] = loan_io_inst_GPIO_OE_bus[35];
assign loanio_gpio_loanio1_oe[7] = loan_io_inst_GPIO_OE_bus[36];
assign loanio_gpio_loanio1_oe[8] = loan_io_inst_GPIO_OE_bus[37];
assign loanio_gpio_loanio1_oe[9] = loan_io_inst_GPIO_OE_bus[38];
assign loanio_gpio_loanio1_oe[10] = loan_io_inst_GPIO_OE_bus[39];
assign loanio_gpio_loanio1_oe[11] = loan_io_inst_GPIO_OE_bus[40];
assign loanio_gpio_loanio1_oe[12] = loan_io_inst_GPIO_OE_bus[41];
assign loanio_gpio_loanio1_oe[13] = loan_io_inst_GPIO_OE_bus[42];
assign loanio_gpio_loanio1_oe[14] = loan_io_inst_GPIO_OE_bus[43];
assign loanio_gpio_loanio1_oe[15] = loan_io_inst_GPIO_OE_bus[44];
assign loanio_gpio_loanio1_oe[16] = loan_io_inst_GPIO_OE_bus[45];
assign loanio_gpio_loanio1_oe[17] = loan_io_inst_GPIO_OE_bus[46];
assign loanio_gpio_loanio1_oe[18] = loan_io_inst_GPIO_OE_bus[47];
assign loanio_gpio_loanio1_oe[19] = loan_io_inst_GPIO_OE_bus[48];
assign loanio_gpio_loanio1_oe[20] = loan_io_inst_GPIO_OE_bus[49];
assign loanio_gpio_loanio1_oe[21] = loan_io_inst_GPIO_OE_bus[50];
assign loanio_gpio_loanio1_oe[22] = loan_io_inst_GPIO_OE_bus[51];
assign loanio_gpio_loanio1_oe[23] = loan_io_inst_GPIO_OE_bus[52];
assign loanio_gpio_loanio1_oe[24] = loan_io_inst_GPIO_OE_bus[53];
assign loanio_gpio_loanio1_oe[25] = loan_io_inst_GPIO_OE_bus[54];
assign loanio_gpio_loanio1_oe[26] = loan_io_inst_GPIO_OE_bus[55];
assign loanio_gpio_loanio1_oe[27] = loan_io_inst_GPIO_OE_bus[56];
assign loanio_gpio_loanio1_oe[28] = loan_io_inst_GPIO_OE_bus[57];
assign loanio_gpio_loanio2_oe[0] = loan_io_inst_GPIO_OE_bus[58];
assign loanio_gpio_loanio2_oe[1] = loan_io_inst_GPIO_OE_bus[59];
assign loanio_gpio_loanio2_oe[2] = loan_io_inst_GPIO_OE_bus[60];
assign loanio_gpio_loanio2_oe[3] = loan_io_inst_GPIO_OE_bus[61];
assign loanio_gpio_loanio2_oe[4] = loan_io_inst_GPIO_OE_bus[62];
assign loanio_gpio_loanio2_oe[5] = loan_io_inst_GPIO_OE_bus[63];
assign loanio_gpio_loanio2_oe[6] = loan_io_inst_GPIO_OE_bus[64];
assign loanio_gpio_loanio2_oe[7] = loan_io_inst_GPIO_OE_bus[65];
assign loanio_gpio_loanio2_oe[8] = loan_io_inst_GPIO_OE_bus[66];

assign loanio_gpio_loanio0_o[0] = loan_io_inst_GPIO_OUT_bus[0];
assign loanio_gpio_loanio0_o[1] = loan_io_inst_GPIO_OUT_bus[1];
assign loanio_gpio_loanio0_o[2] = loan_io_inst_GPIO_OUT_bus[2];
assign loanio_gpio_loanio0_o[3] = loan_io_inst_GPIO_OUT_bus[3];
assign loanio_gpio_loanio0_o[4] = loan_io_inst_GPIO_OUT_bus[4];
assign loanio_gpio_loanio0_o[5] = loan_io_inst_GPIO_OUT_bus[5];
assign loanio_gpio_loanio0_o[6] = loan_io_inst_GPIO_OUT_bus[6];
assign loanio_gpio_loanio0_o[7] = loan_io_inst_GPIO_OUT_bus[7];
assign loanio_gpio_loanio0_o[8] = loan_io_inst_GPIO_OUT_bus[8];
assign loanio_gpio_loanio0_o[9] = loan_io_inst_GPIO_OUT_bus[9];
assign loanio_gpio_loanio0_o[10] = loan_io_inst_GPIO_OUT_bus[10];
assign loanio_gpio_loanio0_o[11] = loan_io_inst_GPIO_OUT_bus[11];
assign loanio_gpio_loanio0_o[12] = loan_io_inst_GPIO_OUT_bus[12];
assign loanio_gpio_loanio0_o[13] = loan_io_inst_GPIO_OUT_bus[13];
assign loanio_gpio_loanio0_o[14] = loan_io_inst_GPIO_OUT_bus[14];
assign loanio_gpio_loanio0_o[15] = loan_io_inst_GPIO_OUT_bus[15];
assign loanio_gpio_loanio0_o[16] = loan_io_inst_GPIO_OUT_bus[16];
assign loanio_gpio_loanio0_o[17] = loan_io_inst_GPIO_OUT_bus[17];
assign loanio_gpio_loanio0_o[18] = loan_io_inst_GPIO_OUT_bus[18];
assign loanio_gpio_loanio0_o[19] = loan_io_inst_GPIO_OUT_bus[19];
assign loanio_gpio_loanio0_o[20] = loan_io_inst_GPIO_OUT_bus[20];
assign loanio_gpio_loanio0_o[21] = loan_io_inst_GPIO_OUT_bus[21];
assign loanio_gpio_loanio0_o[22] = loan_io_inst_GPIO_OUT_bus[22];
assign loanio_gpio_loanio0_o[23] = loan_io_inst_GPIO_OUT_bus[23];
assign loanio_gpio_loanio0_o[24] = loan_io_inst_GPIO_OUT_bus[24];
assign loanio_gpio_loanio0_o[25] = loan_io_inst_GPIO_OUT_bus[25];
assign loanio_gpio_loanio0_o[26] = loan_io_inst_GPIO_OUT_bus[26];
assign loanio_gpio_loanio0_o[27] = loan_io_inst_GPIO_OUT_bus[27];
assign loanio_gpio_loanio0_o[28] = loan_io_inst_GPIO_OUT_bus[28];
assign loanio_gpio_loanio1_o[0] = loan_io_inst_GPIO_OUT_bus[29];
assign loanio_gpio_loanio1_o[1] = loan_io_inst_GPIO_OUT_bus[30];
assign loanio_gpio_loanio1_o[2] = loan_io_inst_GPIO_OUT_bus[31];
assign loanio_gpio_loanio1_o[3] = loan_io_inst_GPIO_OUT_bus[32];
assign loanio_gpio_loanio1_o[4] = loan_io_inst_GPIO_OUT_bus[33];
assign loanio_gpio_loanio1_o[5] = loan_io_inst_GPIO_OUT_bus[34];
assign loanio_gpio_loanio1_o[6] = loan_io_inst_GPIO_OUT_bus[35];
assign loanio_gpio_loanio1_o[7] = loan_io_inst_GPIO_OUT_bus[36];
assign loanio_gpio_loanio1_o[8] = loan_io_inst_GPIO_OUT_bus[37];
assign loanio_gpio_loanio1_o[9] = loan_io_inst_GPIO_OUT_bus[38];
assign loanio_gpio_loanio1_o[10] = loan_io_inst_GPIO_OUT_bus[39];
assign loanio_gpio_loanio1_o[11] = loan_io_inst_GPIO_OUT_bus[40];
assign loanio_gpio_loanio1_o[12] = loan_io_inst_GPIO_OUT_bus[41];
assign loanio_gpio_loanio1_o[13] = loan_io_inst_GPIO_OUT_bus[42];
assign loanio_gpio_loanio1_o[14] = loan_io_inst_GPIO_OUT_bus[43];
assign loanio_gpio_loanio1_o[15] = loan_io_inst_GPIO_OUT_bus[44];
assign loanio_gpio_loanio1_o[16] = loan_io_inst_GPIO_OUT_bus[45];
assign loanio_gpio_loanio1_o[17] = loan_io_inst_GPIO_OUT_bus[46];
assign loanio_gpio_loanio1_o[18] = loan_io_inst_GPIO_OUT_bus[47];
assign loanio_gpio_loanio1_o[19] = loan_io_inst_GPIO_OUT_bus[48];
assign loanio_gpio_loanio1_o[20] = loan_io_inst_GPIO_OUT_bus[49];
assign loanio_gpio_loanio1_o[21] = loan_io_inst_GPIO_OUT_bus[50];
assign loanio_gpio_loanio1_o[22] = loan_io_inst_GPIO_OUT_bus[51];
assign loanio_gpio_loanio1_o[23] = loan_io_inst_GPIO_OUT_bus[52];
assign loanio_gpio_loanio1_o[24] = loan_io_inst_GPIO_OUT_bus[53];
assign loanio_gpio_loanio1_o[25] = loan_io_inst_GPIO_OUT_bus[54];
assign loanio_gpio_loanio1_o[26] = loan_io_inst_GPIO_OUT_bus[55];
assign loanio_gpio_loanio1_o[27] = loan_io_inst_GPIO_OUT_bus[56];
assign loanio_gpio_loanio1_o[28] = loan_io_inst_GPIO_OUT_bus[57];
assign loanio_gpio_loanio2_o[0] = loan_io_inst_GPIO_OUT_bus[58];
assign loanio_gpio_loanio2_o[1] = loan_io_inst_GPIO_OUT_bus[59];
assign loanio_gpio_loanio2_o[2] = loan_io_inst_GPIO_OUT_bus[60];
assign loanio_gpio_loanio2_o[3] = loan_io_inst_GPIO_OUT_bus[61];
assign loanio_gpio_loanio2_o[4] = loan_io_inst_GPIO_OUT_bus[62];
assign loanio_gpio_loanio2_o[5] = loan_io_inst_GPIO_OUT_bus[63];
assign loanio_gpio_loanio2_o[6] = loan_io_inst_GPIO_OUT_bus[64];
assign loanio_gpio_loanio2_o[7] = loan_io_inst_GPIO_OUT_bus[65];
assign loanio_gpio_loanio2_o[8] = loan_io_inst_GPIO_OUT_bus[66];

assign h2f_loan_in[0] = loan_io_inst_LOANIO_IN_bus[0];
assign h2f_loan_in[1] = loan_io_inst_LOANIO_IN_bus[1];
assign h2f_loan_in[2] = loan_io_inst_LOANIO_IN_bus[2];
assign h2f_loan_in[3] = loan_io_inst_LOANIO_IN_bus[3];
assign h2f_loan_in[4] = loan_io_inst_LOANIO_IN_bus[4];
assign h2f_loan_in[5] = loan_io_inst_LOANIO_IN_bus[5];
assign h2f_loan_in[6] = loan_io_inst_LOANIO_IN_bus[6];
assign h2f_loan_in[7] = loan_io_inst_LOANIO_IN_bus[7];
assign h2f_loan_in[8] = loan_io_inst_LOANIO_IN_bus[8];
assign h2f_loan_in[9] = loan_io_inst_LOANIO_IN_bus[9];
assign h2f_loan_in[10] = loan_io_inst_LOANIO_IN_bus[10];
assign h2f_loan_in[11] = loan_io_inst_LOANIO_IN_bus[11];
assign h2f_loan_in[12] = loan_io_inst_LOANIO_IN_bus[12];
assign h2f_loan_in[13] = loan_io_inst_LOANIO_IN_bus[13];
assign h2f_loan_in[14] = loan_io_inst_LOANIO_IN_bus[14];
assign h2f_loan_in[15] = loan_io_inst_LOANIO_IN_bus[15];
assign h2f_loan_in[16] = loan_io_inst_LOANIO_IN_bus[16];
assign h2f_loan_in[17] = loan_io_inst_LOANIO_IN_bus[17];
assign h2f_loan_in[18] = loan_io_inst_LOANIO_IN_bus[18];
assign h2f_loan_in[19] = loan_io_inst_LOANIO_IN_bus[19];
assign h2f_loan_in[20] = loan_io_inst_LOANIO_IN_bus[20];
assign h2f_loan_in[21] = loan_io_inst_LOANIO_IN_bus[21];
assign h2f_loan_in[22] = loan_io_inst_LOANIO_IN_bus[22];
assign h2f_loan_in[23] = loan_io_inst_LOANIO_IN_bus[23];
assign h2f_loan_in[24] = loan_io_inst_LOANIO_IN_bus[24];
assign h2f_loan_in[25] = loan_io_inst_LOANIO_IN_bus[25];
assign h2f_loan_in[26] = loan_io_inst_LOANIO_IN_bus[26];
assign h2f_loan_in[27] = loan_io_inst_LOANIO_IN_bus[27];
assign h2f_loan_in[28] = loan_io_inst_LOANIO_IN_bus[28];
assign h2f_loan_in[29] = loan_io_inst_LOANIO_IN_bus[29];
assign h2f_loan_in[30] = loan_io_inst_LOANIO_IN_bus[30];
assign h2f_loan_in[31] = loan_io_inst_LOANIO_IN_bus[31];
assign h2f_loan_in[32] = loan_io_inst_LOANIO_IN_bus[32];
assign h2f_loan_in[33] = loan_io_inst_LOANIO_IN_bus[33];
assign h2f_loan_in[34] = loan_io_inst_LOANIO_IN_bus[34];
assign h2f_loan_in[35] = loan_io_inst_LOANIO_IN_bus[35];
assign h2f_loan_in[36] = loan_io_inst_LOANIO_IN_bus[36];
assign h2f_loan_in[37] = loan_io_inst_LOANIO_IN_bus[37];
assign h2f_loan_in[38] = loan_io_inst_LOANIO_IN_bus[38];
assign h2f_loan_in[39] = loan_io_inst_LOANIO_IN_bus[39];
assign h2f_loan_in[40] = loan_io_inst_LOANIO_IN_bus[40];
assign h2f_loan_in[41] = loan_io_inst_LOANIO_IN_bus[41];
assign h2f_loan_in[42] = loan_io_inst_LOANIO_IN_bus[42];
assign h2f_loan_in[43] = loan_io_inst_LOANIO_IN_bus[43];
assign h2f_loan_in[44] = loan_io_inst_LOANIO_IN_bus[44];
assign h2f_loan_in[45] = loan_io_inst_LOANIO_IN_bus[45];
assign h2f_loan_in[46] = loan_io_inst_LOANIO_IN_bus[46];
assign h2f_loan_in[47] = loan_io_inst_LOANIO_IN_bus[47];
assign h2f_loan_in[48] = loan_io_inst_LOANIO_IN_bus[48];
assign h2f_loan_in[49] = loan_io_inst_LOANIO_IN_bus[49];
assign h2f_loan_in[50] = loan_io_inst_LOANIO_IN_bus[50];
assign h2f_loan_in[51] = loan_io_inst_LOANIO_IN_bus[51];
assign h2f_loan_in[52] = loan_io_inst_LOANIO_IN_bus[52];
assign h2f_loan_in[53] = loan_io_inst_LOANIO_IN_bus[53];
assign h2f_loan_in[54] = loan_io_inst_LOANIO_IN_bus[54];
assign h2f_loan_in[55] = loan_io_inst_LOANIO_IN_bus[55];
assign h2f_loan_in[56] = loan_io_inst_LOANIO_IN_bus[56];
assign h2f_loan_in[57] = loan_io_inst_LOANIO_IN_bus[57];
assign h2f_loan_in[58] = loan_io_inst_LOANIO_IN_bus[58];
assign h2f_loan_in[59] = loan_io_inst_LOANIO_IN_bus[59];
assign h2f_loan_in[60] = loan_io_inst_LOANIO_IN_bus[60];
assign h2f_loan_in[61] = loan_io_inst_LOANIO_IN_bus[61];
assign h2f_loan_in[62] = loan_io_inst_LOANIO_IN_bus[62];
assign h2f_loan_in[63] = loan_io_inst_LOANIO_IN_bus[63];
assign h2f_loan_in[64] = loan_io_inst_LOANIO_IN_bus[64];
assign h2f_loan_in[65] = loan_io_inst_LOANIO_IN_bus[65];
assign h2f_loan_in[66] = loan_io_inst_LOANIO_IN_bus[66];

assign h2f_lw_ARADDR[0] = hps2fpga_light_weight_ARADDR_bus[0];
assign h2f_lw_ARADDR[1] = hps2fpga_light_weight_ARADDR_bus[1];
assign h2f_lw_ARADDR[2] = hps2fpga_light_weight_ARADDR_bus[2];
assign h2f_lw_ARADDR[3] = hps2fpga_light_weight_ARADDR_bus[3];
assign h2f_lw_ARADDR[4] = hps2fpga_light_weight_ARADDR_bus[4];
assign h2f_lw_ARADDR[5] = hps2fpga_light_weight_ARADDR_bus[5];
assign h2f_lw_ARADDR[6] = hps2fpga_light_weight_ARADDR_bus[6];
assign h2f_lw_ARADDR[7] = hps2fpga_light_weight_ARADDR_bus[7];
assign h2f_lw_ARADDR[8] = hps2fpga_light_weight_ARADDR_bus[8];
assign h2f_lw_ARADDR[9] = hps2fpga_light_weight_ARADDR_bus[9];
assign h2f_lw_ARADDR[10] = hps2fpga_light_weight_ARADDR_bus[10];
assign h2f_lw_ARADDR[11] = hps2fpga_light_weight_ARADDR_bus[11];
assign h2f_lw_ARADDR[12] = hps2fpga_light_weight_ARADDR_bus[12];
assign h2f_lw_ARADDR[13] = hps2fpga_light_weight_ARADDR_bus[13];
assign h2f_lw_ARADDR[14] = hps2fpga_light_weight_ARADDR_bus[14];
assign \h2f_lw_ARADDR[15]  = hps2fpga_light_weight_ARADDR_bus[15];
assign \h2f_lw_ARADDR[16]  = hps2fpga_light_weight_ARADDR_bus[16];
assign \h2f_lw_ARADDR[17]  = hps2fpga_light_weight_ARADDR_bus[17];
assign \h2f_lw_ARADDR[18]  = hps2fpga_light_weight_ARADDR_bus[18];
assign \h2f_lw_ARADDR[19]  = hps2fpga_light_weight_ARADDR_bus[19];
assign \h2f_lw_ARADDR[20]  = hps2fpga_light_weight_ARADDR_bus[20];

assign h2f_lw_ARBURST[0] = hps2fpga_light_weight_ARBURST_bus[0];
assign h2f_lw_ARBURST[1] = hps2fpga_light_weight_ARBURST_bus[1];

assign h2f_lw_ARID[0] = hps2fpga_light_weight_ARID_bus[0];
assign h2f_lw_ARID[1] = hps2fpga_light_weight_ARID_bus[1];
assign h2f_lw_ARID[2] = hps2fpga_light_weight_ARID_bus[2];
assign h2f_lw_ARID[3] = hps2fpga_light_weight_ARID_bus[3];
assign h2f_lw_ARID[4] = hps2fpga_light_weight_ARID_bus[4];
assign h2f_lw_ARID[5] = hps2fpga_light_weight_ARID_bus[5];
assign h2f_lw_ARID[6] = hps2fpga_light_weight_ARID_bus[6];
assign h2f_lw_ARID[7] = hps2fpga_light_weight_ARID_bus[7];
assign h2f_lw_ARID[8] = hps2fpga_light_weight_ARID_bus[8];
assign h2f_lw_ARID[9] = hps2fpga_light_weight_ARID_bus[9];
assign h2f_lw_ARID[10] = hps2fpga_light_weight_ARID_bus[10];
assign h2f_lw_ARID[11] = hps2fpga_light_weight_ARID_bus[11];

assign h2f_lw_ARLEN[0] = hps2fpga_light_weight_ARLEN_bus[0];
assign h2f_lw_ARLEN[1] = hps2fpga_light_weight_ARLEN_bus[1];
assign h2f_lw_ARLEN[2] = hps2fpga_light_weight_ARLEN_bus[2];
assign h2f_lw_ARLEN[3] = hps2fpga_light_weight_ARLEN_bus[3];

assign h2f_lw_ARSIZE[0] = hps2fpga_light_weight_ARSIZE_bus[0];
assign h2f_lw_ARSIZE[1] = hps2fpga_light_weight_ARSIZE_bus[1];
assign h2f_lw_ARSIZE[2] = hps2fpga_light_weight_ARSIZE_bus[2];

assign h2f_lw_AWADDR[0] = hps2fpga_light_weight_AWADDR_bus[0];
assign h2f_lw_AWADDR[1] = hps2fpga_light_weight_AWADDR_bus[1];
assign h2f_lw_AWADDR[2] = hps2fpga_light_weight_AWADDR_bus[2];
assign h2f_lw_AWADDR[3] = hps2fpga_light_weight_AWADDR_bus[3];
assign h2f_lw_AWADDR[4] = hps2fpga_light_weight_AWADDR_bus[4];
assign h2f_lw_AWADDR[5] = hps2fpga_light_weight_AWADDR_bus[5];
assign h2f_lw_AWADDR[6] = hps2fpga_light_weight_AWADDR_bus[6];
assign h2f_lw_AWADDR[7] = hps2fpga_light_weight_AWADDR_bus[7];
assign h2f_lw_AWADDR[8] = hps2fpga_light_weight_AWADDR_bus[8];
assign h2f_lw_AWADDR[9] = hps2fpga_light_weight_AWADDR_bus[9];
assign h2f_lw_AWADDR[10] = hps2fpga_light_weight_AWADDR_bus[10];
assign h2f_lw_AWADDR[11] = hps2fpga_light_weight_AWADDR_bus[11];
assign h2f_lw_AWADDR[12] = hps2fpga_light_weight_AWADDR_bus[12];
assign h2f_lw_AWADDR[13] = hps2fpga_light_weight_AWADDR_bus[13];
assign h2f_lw_AWADDR[14] = hps2fpga_light_weight_AWADDR_bus[14];

assign h2f_lw_AWBURST[0] = hps2fpga_light_weight_AWBURST_bus[0];
assign h2f_lw_AWBURST[1] = hps2fpga_light_weight_AWBURST_bus[1];

assign h2f_lw_AWID[0] = hps2fpga_light_weight_AWID_bus[0];
assign h2f_lw_AWID[1] = hps2fpga_light_weight_AWID_bus[1];
assign h2f_lw_AWID[2] = hps2fpga_light_weight_AWID_bus[2];
assign h2f_lw_AWID[3] = hps2fpga_light_weight_AWID_bus[3];
assign h2f_lw_AWID[4] = hps2fpga_light_weight_AWID_bus[4];
assign h2f_lw_AWID[5] = hps2fpga_light_weight_AWID_bus[5];
assign h2f_lw_AWID[6] = hps2fpga_light_weight_AWID_bus[6];
assign h2f_lw_AWID[7] = hps2fpga_light_weight_AWID_bus[7];
assign h2f_lw_AWID[8] = hps2fpga_light_weight_AWID_bus[8];
assign h2f_lw_AWID[9] = hps2fpga_light_weight_AWID_bus[9];
assign h2f_lw_AWID[10] = hps2fpga_light_weight_AWID_bus[10];
assign h2f_lw_AWID[11] = hps2fpga_light_weight_AWID_bus[11];

assign h2f_lw_AWLEN[0] = hps2fpga_light_weight_AWLEN_bus[0];
assign h2f_lw_AWLEN[1] = hps2fpga_light_weight_AWLEN_bus[1];
assign h2f_lw_AWLEN[2] = hps2fpga_light_weight_AWLEN_bus[2];
assign h2f_lw_AWLEN[3] = hps2fpga_light_weight_AWLEN_bus[3];

assign h2f_lw_AWSIZE[0] = hps2fpga_light_weight_AWSIZE_bus[0];
assign h2f_lw_AWSIZE[1] = hps2fpga_light_weight_AWSIZE_bus[1];
assign h2f_lw_AWSIZE[2] = hps2fpga_light_weight_AWSIZE_bus[2];

assign h2f_lw_WDATA[0] = hps2fpga_light_weight_WDATA_bus[0];
assign h2f_lw_WDATA[1] = hps2fpga_light_weight_WDATA_bus[1];
assign h2f_lw_WDATA[2] = hps2fpga_light_weight_WDATA_bus[2];
assign h2f_lw_WDATA[3] = hps2fpga_light_weight_WDATA_bus[3];
assign h2f_lw_WDATA[4] = hps2fpga_light_weight_WDATA_bus[4];
assign h2f_lw_WDATA[5] = hps2fpga_light_weight_WDATA_bus[5];
assign h2f_lw_WDATA[6] = hps2fpga_light_weight_WDATA_bus[6];
assign h2f_lw_WDATA[7] = hps2fpga_light_weight_WDATA_bus[7];
assign h2f_lw_WDATA[8] = hps2fpga_light_weight_WDATA_bus[8];
assign h2f_lw_WDATA[9] = hps2fpga_light_weight_WDATA_bus[9];
assign h2f_lw_WDATA[10] = hps2fpga_light_weight_WDATA_bus[10];
assign h2f_lw_WDATA[11] = hps2fpga_light_weight_WDATA_bus[11];
assign h2f_lw_WDATA[12] = hps2fpga_light_weight_WDATA_bus[12];
assign h2f_lw_WDATA[13] = hps2fpga_light_weight_WDATA_bus[13];
assign h2f_lw_WDATA[14] = hps2fpga_light_weight_WDATA_bus[14];
assign h2f_lw_WDATA[15] = hps2fpga_light_weight_WDATA_bus[15];
assign h2f_lw_WDATA[16] = hps2fpga_light_weight_WDATA_bus[16];
assign h2f_lw_WDATA[17] = hps2fpga_light_weight_WDATA_bus[17];
assign h2f_lw_WDATA[18] = hps2fpga_light_weight_WDATA_bus[18];
assign h2f_lw_WDATA[19] = hps2fpga_light_weight_WDATA_bus[19];
assign h2f_lw_WDATA[20] = hps2fpga_light_weight_WDATA_bus[20];
assign h2f_lw_WDATA[21] = hps2fpga_light_weight_WDATA_bus[21];
assign h2f_lw_WDATA[22] = hps2fpga_light_weight_WDATA_bus[22];
assign h2f_lw_WDATA[23] = hps2fpga_light_weight_WDATA_bus[23];
assign h2f_lw_WDATA[24] = hps2fpga_light_weight_WDATA_bus[24];
assign h2f_lw_WDATA[25] = hps2fpga_light_weight_WDATA_bus[25];
assign h2f_lw_WDATA[26] = hps2fpga_light_weight_WDATA_bus[26];
assign h2f_lw_WDATA[27] = hps2fpga_light_weight_WDATA_bus[27];
assign h2f_lw_WDATA[28] = hps2fpga_light_weight_WDATA_bus[28];
assign h2f_lw_WDATA[29] = hps2fpga_light_weight_WDATA_bus[29];
assign h2f_lw_WDATA[30] = hps2fpga_light_weight_WDATA_bus[30];
assign h2f_lw_WDATA[31] = hps2fpga_light_weight_WDATA_bus[31];

assign h2f_lw_WSTRB[0] = hps2fpga_light_weight_WSTRB_bus[0];
assign h2f_lw_WSTRB[1] = hps2fpga_light_weight_WSTRB_bus[1];
assign h2f_lw_WSTRB[2] = hps2fpga_light_weight_WSTRB_bus[2];
assign h2f_lw_WSTRB[3] = hps2fpga_light_weight_WSTRB_bus[3];

cyclonev_hps_interface_loan_io loan_io_inst(
	.gpio_in({gnd,gnd,gnd,gnd,loanio_gpio_loanio2_i[8],loanio_gpio_loanio2_i[7],loanio_gpio_loanio2_i[6],loanio_gpio_loanio2_i[5],loanio_gpio_loanio2_i[4],loanio_gpio_loanio2_i[3],loanio_gpio_loanio2_i[2],loanio_gpio_loanio2_i[1],loanio_gpio_loanio2_i[0],loanio_gpio_loanio1_i[28],loanio_gpio_loanio1_i[27],
loanio_gpio_loanio1_i[26],loanio_gpio_loanio1_i[25],loanio_gpio_loanio1_i[24],loanio_gpio_loanio1_i[23],loanio_gpio_loanio1_i[22],loanio_gpio_loanio1_i[21],loanio_gpio_loanio1_i[20],loanio_gpio_loanio1_i[19],loanio_gpio_loanio1_i[18],loanio_gpio_loanio1_i[17],loanio_gpio_loanio1_i[16],loanio_gpio_loanio1_i[15],
loanio_gpio_loanio1_i[14],loanio_gpio_loanio1_i[13],loanio_gpio_loanio1_i[12],loanio_gpio_loanio1_i[11],loanio_gpio_loanio1_i[10],loanio_gpio_loanio1_i[9],loanio_gpio_loanio1_i[8],loanio_gpio_loanio1_i[7],loanio_gpio_loanio1_i[6],loanio_gpio_loanio1_i[5],loanio_gpio_loanio1_i[4],loanio_gpio_loanio1_i[3],
loanio_gpio_loanio1_i[2],loanio_gpio_loanio1_i[1],loanio_gpio_loanio1_i[0],loanio_gpio_loanio0_i[28],loanio_gpio_loanio0_i[27],loanio_gpio_loanio0_i[26],loanio_gpio_loanio0_i[25],loanio_gpio_loanio0_i[24],loanio_gpio_loanio0_i[23],loanio_gpio_loanio0_i[22],loanio_gpio_loanio0_i[21],loanio_gpio_loanio0_i[20],
loanio_gpio_loanio0_i[19],loanio_gpio_loanio0_i[18],loanio_gpio_loanio0_i[17],loanio_gpio_loanio0_i[16],loanio_gpio_loanio0_i[15],loanio_gpio_loanio0_i[14],loanio_gpio_loanio0_i[13],loanio_gpio_loanio0_i[12],loanio_gpio_loanio0_i[11],loanio_gpio_loanio0_i[10],loanio_gpio_loanio0_i[9],loanio_gpio_loanio0_i[8],
loanio_gpio_loanio0_i[7],loanio_gpio_loanio0_i[6],loanio_gpio_loanio0_i[5],loanio_gpio_loanio0_i[4],loanio_gpio_loanio0_i[3],loanio_gpio_loanio0_i[2],loanio_gpio_loanio0_i[1],loanio_gpio_loanio0_i[0]}),
	.loanio_oe({gnd,gnd,gnd,gnd,h2f_loan_oe[66],h2f_loan_oe[65],h2f_loan_oe[64],h2f_loan_oe[63],h2f_loan_oe[62],h2f_loan_oe[61],h2f_loan_oe[60],h2f_loan_oe[59],h2f_loan_oe[58],h2f_loan_oe[57],h2f_loan_oe[56],h2f_loan_oe[55],h2f_loan_oe[54],h2f_loan_oe[53],h2f_loan_oe[52],h2f_loan_oe[51],h2f_loan_oe[50],h2f_loan_oe[49],h2f_loan_oe[48],h2f_loan_oe[47],h2f_loan_oe[46],h2f_loan_oe[45],
h2f_loan_oe[44],h2f_loan_oe[43],h2f_loan_oe[42],h2f_loan_oe[41],h2f_loan_oe[40],h2f_loan_oe[39],h2f_loan_oe[38],h2f_loan_oe[37],h2f_loan_oe[36],h2f_loan_oe[35],h2f_loan_oe[34],h2f_loan_oe[33],h2f_loan_oe[32],h2f_loan_oe[31],h2f_loan_oe[30],h2f_loan_oe[29],h2f_loan_oe[28],h2f_loan_oe[27],h2f_loan_oe[26],h2f_loan_oe[25],h2f_loan_oe[24],h2f_loan_oe[23],h2f_loan_oe[22],
h2f_loan_oe[21],h2f_loan_oe[20],h2f_loan_oe[19],h2f_loan_oe[18],h2f_loan_oe[17],h2f_loan_oe[16],h2f_loan_oe[15],h2f_loan_oe[14],h2f_loan_oe[13],h2f_loan_oe[12],h2f_loan_oe[11],h2f_loan_oe[10],h2f_loan_oe[9],h2f_loan_oe[8],h2f_loan_oe[7],h2f_loan_oe[6],h2f_loan_oe[5],h2f_loan_oe[4],h2f_loan_oe[3],h2f_loan_oe[2],h2f_loan_oe[1],h2f_loan_oe[0]}),
	.loanio_out({gnd,gnd,gnd,gnd,h2f_loan_out[66],h2f_loan_out[65],h2f_loan_out[64],h2f_loan_out[63],h2f_loan_out[62],h2f_loan_out[61],h2f_loan_out[60],h2f_loan_out[59],h2f_loan_out[58],h2f_loan_out[57],h2f_loan_out[56],h2f_loan_out[55],h2f_loan_out[54],h2f_loan_out[53],h2f_loan_out[52],h2f_loan_out[51],h2f_loan_out[50],h2f_loan_out[49],h2f_loan_out[48],h2f_loan_out[47],
h2f_loan_out[46],h2f_loan_out[45],h2f_loan_out[44],h2f_loan_out[43],h2f_loan_out[42],h2f_loan_out[41],h2f_loan_out[40],h2f_loan_out[39],h2f_loan_out[38],h2f_loan_out[37],h2f_loan_out[36],h2f_loan_out[35],h2f_loan_out[34],h2f_loan_out[33],h2f_loan_out[32],h2f_loan_out[31],h2f_loan_out[30],h2f_loan_out[29],h2f_loan_out[28],h2f_loan_out[27],h2f_loan_out[26],
h2f_loan_out[25],h2f_loan_out[24],h2f_loan_out[23],h2f_loan_out[22],h2f_loan_out[21],h2f_loan_out[20],h2f_loan_out[19],h2f_loan_out[18],h2f_loan_out[17],h2f_loan_out[16],h2f_loan_out[15],h2f_loan_out[14],h2f_loan_out[13],h2f_loan_out[12],h2f_loan_out[11],h2f_loan_out[10],h2f_loan_out[9],h2f_loan_out[8],h2f_loan_out[7],h2f_loan_out[6],h2f_loan_out[5],
h2f_loan_out[4],h2f_loan_out[3],h2f_loan_out[2],h2f_loan_out[1],h2f_loan_out[0]}),
	.fake_dout(\loan_io_inst~fake_dout ),
	.gpio_oe(loan_io_inst_GPIO_OE_bus),
	.gpio_out(loan_io_inst_GPIO_OUT_bus),
	.input_only(),
	.loanio_in(loan_io_inst_LOANIO_IN_bus));

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(vcc),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(\clocks_resets~h2f_cold_rst_n ),
	.h2f_pending_rst_req_n(),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_hps2fpga_light_weight hps2fpga_light_weight(
	.arready(h2f_lw_ARREADY[0]),
	.awready(h2f_lw_AWREADY[0]),
	.bvalid(h2f_lw_BVALID[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(h2f_lw_RLAST[0]),
	.rvalid(h2f_lw_RVALID[0]),
	.wready(h2f_lw_WREADY[0]),
	.bid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.bresp({gnd,gnd}),
	.rdata({h2f_lw_RDATA[31],h2f_lw_RDATA[30],h2f_lw_RDATA[29],h2f_lw_RDATA[28],h2f_lw_RDATA[27],h2f_lw_RDATA[26],h2f_lw_RDATA[25],h2f_lw_RDATA[24],h2f_lw_RDATA[23],h2f_lw_RDATA[22],h2f_lw_RDATA[21],h2f_lw_RDATA[20],h2f_lw_RDATA[19],h2f_lw_RDATA[18],h2f_lw_RDATA[17],h2f_lw_RDATA[16],h2f_lw_RDATA[15],h2f_lw_RDATA[14],h2f_lw_RDATA[13],h2f_lw_RDATA[12],h2f_lw_RDATA[11],
h2f_lw_RDATA[10],h2f_lw_RDATA[9],h2f_lw_RDATA[8],h2f_lw_RDATA[7],h2f_lw_RDATA[6],h2f_lw_RDATA[5],h2f_lw_RDATA[4],h2f_lw_RDATA[3],h2f_lw_RDATA[2],h2f_lw_RDATA[1],h2f_lw_RDATA[0]}),
	.rid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_lw_ARVALID[0]),
	.awvalid(h2f_lw_AWVALID[0]),
	.bready(h2f_lw_BREADY[0]),
	.rready(h2f_lw_RREADY[0]),
	.wlast(h2f_lw_WLAST[0]),
	.wvalid(h2f_lw_WVALID[0]),
	.araddr(hps2fpga_light_weight_ARADDR_bus),
	.arburst(hps2fpga_light_weight_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_light_weight_ARID_bus),
	.arlen(hps2fpga_light_weight_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_light_weight_ARSIZE_bus),
	.awaddr(hps2fpga_light_weight_AWADDR_bus),
	.awburst(hps2fpga_light_weight_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_light_weight_AWID_bus),
	.awlen(hps2fpga_light_weight_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_light_weight_AWSIZE_bus),
	.wdata(hps2fpga_light_weight_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_light_weight_WSTRB_bus));

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(gnd),
	.awvalid(gnd),
	.bready(gnd),
	.clk(gnd),
	.rready(gnd),
	.wlast(gnd),
	.wvalid(gnd),
	.araddr(32'b00000000000000000000000000000000),
	.arburst(2'b00),
	.arcache(4'b0000),
	.arid(8'b00000000),
	.arlen(4'b0000),
	.arlock(2'b00),
	.arprot(3'b000),
	.arsize(3'b000),
	.aruser(5'b00000),
	.awaddr(32'b00000000000000000000000000000000),
	.awburst(2'b00),
	.awcache(4'b0000),
	.awid(8'b00000000),
	.awlen(4'b0000),
	.awlock(2'b00),
	.awprot(3'b000),
	.awsize(3'b000),
	.awuser(5'b00000),
	.port_size_config({vcc,vcc}),
	.wdata(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wid(8'b00000000),
	.wstrb(16'b0000000000000000),
	.arready(\fpga2hps~arready ),
	.awready(),
	.bvalid(),
	.rlast(),
	.rvalid(),
	.wready(),
	.bid(),
	.bresp(),
	.rdata(),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(gnd),
	.awready(gnd),
	.bvalid(gnd),
	.clk(gnd),
	.rlast(gnd),
	.rvalid(gnd),
	.wready(gnd),
	.bid(12'b000000000000),
	.bresp(2'b00),
	.port_size_config({vcc,vcc}),
	.rdata(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.rid(12'b000000000000),
	.rresp(2'b00),
	.arvalid(),
	.awvalid(),
	.bready(),
	.rready(),
	.wlast(),
	.wvalid(),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(),
	.arcache(),
	.arid(),
	.arlen(),
	.arlock(),
	.arprot(),
	.arsize(),
	.awaddr(),
	.awburst(),
	.awcache(),
	.awid(),
	.awlen(),
	.awlock(),
	.awprot(),
	.awsize(),
	.wdata(),
	.wid(),
	.wstrb());
defparam hps2fpga.data_width = 32;

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(gnd),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(gnd),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(gnd),
	.rd_clk_1(gnd),
	.rd_clk_2(gnd),
	.rd_clk_3(gnd),
	.rd_ready_0(gnd),
	.rd_ready_1(gnd),
	.rd_ready_2(gnd),
	.rd_ready_3(gnd),
	.wr_clk_0(gnd),
	.wr_clk_1(gnd),
	.wr_clk_2(gnd),
	.wr_clk_3(gnd),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(gnd),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_1(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_2(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_3(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.cmd_ready_0(),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(),
	.rd_data_1(),
	.rd_data_2(),
	.rd_data_3(),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

endmodule

module soc_system_soc_system_hps_0_hps_io (
	loanio_gpio_loanio0_oe_0,
	loanio_gpio_loanio0_oe_1,
	loanio_gpio_loanio0_oe_2,
	loanio_gpio_loanio0_oe_3,
	loanio_gpio_loanio0_oe_4,
	loanio_gpio_loanio0_oe_5,
	loanio_gpio_loanio0_oe_6,
	loanio_gpio_loanio0_oe_7,
	loanio_gpio_loanio0_oe_8,
	loanio_gpio_loanio0_oe_9,
	loanio_gpio_loanio0_oe_10,
	loanio_gpio_loanio0_oe_11,
	loanio_gpio_loanio0_oe_12,
	loanio_gpio_loanio0_oe_13,
	loanio_gpio_loanio0_oe_14,
	loanio_gpio_loanio0_oe_15,
	loanio_gpio_loanio0_oe_16,
	loanio_gpio_loanio0_oe_17,
	loanio_gpio_loanio0_oe_18,
	loanio_gpio_loanio0_oe_19,
	loanio_gpio_loanio0_oe_20,
	loanio_gpio_loanio0_oe_21,
	loanio_gpio_loanio0_oe_22,
	loanio_gpio_loanio0_oe_23,
	loanio_gpio_loanio0_oe_24,
	loanio_gpio_loanio0_oe_25,
	loanio_gpio_loanio0_oe_26,
	loanio_gpio_loanio0_oe_27,
	loanio_gpio_loanio0_oe_28,
	loanio_gpio_loanio1_oe_0,
	loanio_gpio_loanio1_oe_1,
	loanio_gpio_loanio1_oe_2,
	loanio_gpio_loanio1_oe_3,
	loanio_gpio_loanio1_oe_4,
	loanio_gpio_loanio1_oe_5,
	loanio_gpio_loanio1_oe_6,
	loanio_gpio_loanio1_oe_7,
	loanio_gpio_loanio1_oe_8,
	loanio_gpio_loanio1_oe_9,
	loanio_gpio_loanio1_oe_10,
	loanio_gpio_loanio1_oe_11,
	loanio_gpio_loanio1_oe_12,
	loanio_gpio_loanio1_oe_13,
	loanio_gpio_loanio1_oe_14,
	loanio_gpio_loanio1_oe_15,
	loanio_gpio_loanio1_oe_16,
	loanio_gpio_loanio1_oe_17,
	loanio_gpio_loanio1_oe_18,
	loanio_gpio_loanio1_oe_19,
	loanio_gpio_loanio1_oe_20,
	loanio_gpio_loanio1_oe_21,
	loanio_gpio_loanio1_oe_22,
	loanio_gpio_loanio1_oe_23,
	loanio_gpio_loanio1_oe_24,
	loanio_gpio_loanio1_oe_25,
	loanio_gpio_loanio1_oe_26,
	loanio_gpio_loanio1_oe_27,
	loanio_gpio_loanio1_oe_28,
	loanio_gpio_loanio2_oe_0,
	loanio_gpio_loanio2_oe_1,
	loanio_gpio_loanio2_oe_2,
	loanio_gpio_loanio2_oe_3,
	loanio_gpio_loanio2_oe_4,
	loanio_gpio_loanio2_oe_5,
	loanio_gpio_loanio2_oe_6,
	loanio_gpio_loanio2_oe_7,
	loanio_gpio_loanio2_oe_8,
	loanio_gpio_loanio0_o_0,
	loanio_gpio_loanio0_o_1,
	loanio_gpio_loanio0_o_2,
	loanio_gpio_loanio0_o_3,
	loanio_gpio_loanio0_o_4,
	loanio_gpio_loanio0_o_5,
	loanio_gpio_loanio0_o_6,
	loanio_gpio_loanio0_o_7,
	loanio_gpio_loanio0_o_8,
	loanio_gpio_loanio0_o_9,
	loanio_gpio_loanio0_o_10,
	loanio_gpio_loanio0_o_11,
	loanio_gpio_loanio0_o_12,
	loanio_gpio_loanio0_o_13,
	loanio_gpio_loanio0_o_14,
	loanio_gpio_loanio0_o_15,
	loanio_gpio_loanio0_o_16,
	loanio_gpio_loanio0_o_17,
	loanio_gpio_loanio0_o_18,
	loanio_gpio_loanio0_o_19,
	loanio_gpio_loanio0_o_20,
	loanio_gpio_loanio0_o_21,
	loanio_gpio_loanio0_o_22,
	loanio_gpio_loanio0_o_23,
	loanio_gpio_loanio0_o_24,
	loanio_gpio_loanio0_o_25,
	loanio_gpio_loanio0_o_26,
	loanio_gpio_loanio0_o_27,
	loanio_gpio_loanio0_o_28,
	loanio_gpio_loanio1_o_0,
	loanio_gpio_loanio1_o_1,
	loanio_gpio_loanio1_o_2,
	loanio_gpio_loanio1_o_3,
	loanio_gpio_loanio1_o_4,
	loanio_gpio_loanio1_o_5,
	loanio_gpio_loanio1_o_6,
	loanio_gpio_loanio1_o_7,
	loanio_gpio_loanio1_o_8,
	loanio_gpio_loanio1_o_9,
	loanio_gpio_loanio1_o_10,
	loanio_gpio_loanio1_o_11,
	loanio_gpio_loanio1_o_12,
	loanio_gpio_loanio1_o_13,
	loanio_gpio_loanio1_o_14,
	loanio_gpio_loanio1_o_15,
	loanio_gpio_loanio1_o_16,
	loanio_gpio_loanio1_o_17,
	loanio_gpio_loanio1_o_18,
	loanio_gpio_loanio1_o_19,
	loanio_gpio_loanio1_o_20,
	loanio_gpio_loanio1_o_21,
	loanio_gpio_loanio1_o_22,
	loanio_gpio_loanio1_o_23,
	loanio_gpio_loanio1_o_24,
	loanio_gpio_loanio1_o_25,
	loanio_gpio_loanio1_o_26,
	loanio_gpio_loanio1_o_27,
	loanio_gpio_loanio1_o_28,
	loanio_gpio_loanio2_o_0,
	loanio_gpio_loanio2_o_1,
	loanio_gpio_loanio2_o_2,
	loanio_gpio_loanio2_o_3,
	loanio_gpio_loanio2_o_4,
	loanio_gpio_loanio2_o_5,
	loanio_gpio_loanio2_o_6,
	loanio_gpio_loanio2_o_7,
	loanio_gpio_loanio2_o_8,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim0_inst,
	spim0_inst1,
	intermediate_36,
	intermediate_37,
	spim1_inst,
	spim1_inst1,
	intermediate_38,
	intermediate_39,
	uart0_inst,
	gpio_inst,
	gpio_inst1,
	gpio_inst2,
	gpio_inst3,
	gpio_inst4,
	gpio_inst5,
	gpio_inst6,
	gpio_inst7,
	gpio_inst8,
	gpio_inst9,
	gpio_inst10,
	gpio_inst11,
	gpio_inst12,
	gpio_inst13,
	gpio_inst14,
	gpio_inst15,
	gpio_inst16,
	gpio_inst17,
	gpio_inst18,
	gpio_inst19,
	gpio_inst20,
	gpio_inst21,
	gpio_inst22,
	gpio_inst23,
	gpio_inst24,
	gpio_inst25,
	gpio_inst26,
	gpio_inst27,
	gpio_inst28,
	gpio_inst29,
	gpio_inst30,
	gpio_inst31,
	gpio_inst32,
	gpio_inst33,
	gpio_inst34,
	gpio_inst35,
	gpio_inst36,
	gpio_inst37,
	gpio_inst38,
	gpio_inst39,
	gpio_inst40,
	gpio_inst41,
	gpio_inst42,
	gpio_inst43,
	gpio_inst44,
	gpio_inst45,
	gpio_inst46,
	gpio_inst47,
	gpio_inst48,
	gpio_inst49,
	gpio_inst50,
	gpio_inst51,
	gpio_inst52,
	gpio_inst53,
	gpio_inst54,
	gpio_inst55,
	gpio_inst56,
	gpio_inst57,
	gpio_inst58,
	gpio_inst59,
	gpio_inst60,
	gpio_inst61,
	gpio_inst62,
	gpio_inst63,
	gpio_inst64,
	gpio_inst65,
	gpio_inst66,
	intermediate_50,
	intermediate_40,
	intermediate_51,
	intermediate_41,
	intermediate_42,
	intermediate_52,
	intermediate_44,
	intermediate_54,
	intermediate_56,
	intermediate_58,
	intermediate_60,
	intermediate_62,
	intermediate_64,
	intermediate_43,
	intermediate_53,
	intermediate_45,
	intermediate_55,
	intermediate_57,
	intermediate_59,
	intermediate_61,
	intermediate_63,
	intermediate_65,
	intermediate_46,
	intermediate_48,
	intermediate_47,
	intermediate_49,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_gpio_inst_GPIO62_0,
	hps_io_gpio_inst_LOANIO00_0,
	hps_io_gpio_inst_LOANIO41_0,
	hps_io_gpio_inst_LOANIO51_0,
	hps_io_gpio_inst_LOANIO52_0,
	hps_io_gpio_inst_LOANIO53_0,
	hps_io_gpio_inst_LOANIO54_0,
	hps_io_gpio_inst_LOANIO55_0,
	hps_io_gpio_inst_LOANIO56_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim0_inst_MISO,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
input 	loanio_gpio_loanio0_oe_0;
input 	loanio_gpio_loanio0_oe_1;
input 	loanio_gpio_loanio0_oe_2;
input 	loanio_gpio_loanio0_oe_3;
input 	loanio_gpio_loanio0_oe_4;
input 	loanio_gpio_loanio0_oe_5;
input 	loanio_gpio_loanio0_oe_6;
input 	loanio_gpio_loanio0_oe_7;
input 	loanio_gpio_loanio0_oe_8;
input 	loanio_gpio_loanio0_oe_9;
input 	loanio_gpio_loanio0_oe_10;
input 	loanio_gpio_loanio0_oe_11;
input 	loanio_gpio_loanio0_oe_12;
input 	loanio_gpio_loanio0_oe_13;
input 	loanio_gpio_loanio0_oe_14;
input 	loanio_gpio_loanio0_oe_15;
input 	loanio_gpio_loanio0_oe_16;
input 	loanio_gpio_loanio0_oe_17;
input 	loanio_gpio_loanio0_oe_18;
input 	loanio_gpio_loanio0_oe_19;
input 	loanio_gpio_loanio0_oe_20;
input 	loanio_gpio_loanio0_oe_21;
input 	loanio_gpio_loanio0_oe_22;
input 	loanio_gpio_loanio0_oe_23;
input 	loanio_gpio_loanio0_oe_24;
input 	loanio_gpio_loanio0_oe_25;
input 	loanio_gpio_loanio0_oe_26;
input 	loanio_gpio_loanio0_oe_27;
input 	loanio_gpio_loanio0_oe_28;
input 	loanio_gpio_loanio1_oe_0;
input 	loanio_gpio_loanio1_oe_1;
input 	loanio_gpio_loanio1_oe_2;
input 	loanio_gpio_loanio1_oe_3;
input 	loanio_gpio_loanio1_oe_4;
input 	loanio_gpio_loanio1_oe_5;
input 	loanio_gpio_loanio1_oe_6;
input 	loanio_gpio_loanio1_oe_7;
input 	loanio_gpio_loanio1_oe_8;
input 	loanio_gpio_loanio1_oe_9;
input 	loanio_gpio_loanio1_oe_10;
input 	loanio_gpio_loanio1_oe_11;
input 	loanio_gpio_loanio1_oe_12;
input 	loanio_gpio_loanio1_oe_13;
input 	loanio_gpio_loanio1_oe_14;
input 	loanio_gpio_loanio1_oe_15;
input 	loanio_gpio_loanio1_oe_16;
input 	loanio_gpio_loanio1_oe_17;
input 	loanio_gpio_loanio1_oe_18;
input 	loanio_gpio_loanio1_oe_19;
input 	loanio_gpio_loanio1_oe_20;
input 	loanio_gpio_loanio1_oe_21;
input 	loanio_gpio_loanio1_oe_22;
input 	loanio_gpio_loanio1_oe_23;
input 	loanio_gpio_loanio1_oe_24;
input 	loanio_gpio_loanio1_oe_25;
input 	loanio_gpio_loanio1_oe_26;
input 	loanio_gpio_loanio1_oe_27;
input 	loanio_gpio_loanio1_oe_28;
input 	loanio_gpio_loanio2_oe_0;
input 	loanio_gpio_loanio2_oe_1;
input 	loanio_gpio_loanio2_oe_2;
input 	loanio_gpio_loanio2_oe_3;
input 	loanio_gpio_loanio2_oe_4;
input 	loanio_gpio_loanio2_oe_5;
input 	loanio_gpio_loanio2_oe_6;
input 	loanio_gpio_loanio2_oe_7;
input 	loanio_gpio_loanio2_oe_8;
input 	loanio_gpio_loanio0_o_0;
input 	loanio_gpio_loanio0_o_1;
input 	loanio_gpio_loanio0_o_2;
input 	loanio_gpio_loanio0_o_3;
input 	loanio_gpio_loanio0_o_4;
input 	loanio_gpio_loanio0_o_5;
input 	loanio_gpio_loanio0_o_6;
input 	loanio_gpio_loanio0_o_7;
input 	loanio_gpio_loanio0_o_8;
input 	loanio_gpio_loanio0_o_9;
input 	loanio_gpio_loanio0_o_10;
input 	loanio_gpio_loanio0_o_11;
input 	loanio_gpio_loanio0_o_12;
input 	loanio_gpio_loanio0_o_13;
input 	loanio_gpio_loanio0_o_14;
input 	loanio_gpio_loanio0_o_15;
input 	loanio_gpio_loanio0_o_16;
input 	loanio_gpio_loanio0_o_17;
input 	loanio_gpio_loanio0_o_18;
input 	loanio_gpio_loanio0_o_19;
input 	loanio_gpio_loanio0_o_20;
input 	loanio_gpio_loanio0_o_21;
input 	loanio_gpio_loanio0_o_22;
input 	loanio_gpio_loanio0_o_23;
input 	loanio_gpio_loanio0_o_24;
input 	loanio_gpio_loanio0_o_25;
input 	loanio_gpio_loanio0_o_26;
input 	loanio_gpio_loanio0_o_27;
input 	loanio_gpio_loanio0_o_28;
input 	loanio_gpio_loanio1_o_0;
input 	loanio_gpio_loanio1_o_1;
input 	loanio_gpio_loanio1_o_2;
input 	loanio_gpio_loanio1_o_3;
input 	loanio_gpio_loanio1_o_4;
input 	loanio_gpio_loanio1_o_5;
input 	loanio_gpio_loanio1_o_6;
input 	loanio_gpio_loanio1_o_7;
input 	loanio_gpio_loanio1_o_8;
input 	loanio_gpio_loanio1_o_9;
input 	loanio_gpio_loanio1_o_10;
input 	loanio_gpio_loanio1_o_11;
input 	loanio_gpio_loanio1_o_12;
input 	loanio_gpio_loanio1_o_13;
input 	loanio_gpio_loanio1_o_14;
input 	loanio_gpio_loanio1_o_15;
input 	loanio_gpio_loanio1_o_16;
input 	loanio_gpio_loanio1_o_17;
input 	loanio_gpio_loanio1_o_18;
input 	loanio_gpio_loanio1_o_19;
input 	loanio_gpio_loanio1_o_20;
input 	loanio_gpio_loanio1_o_21;
input 	loanio_gpio_loanio1_o_22;
input 	loanio_gpio_loanio1_o_23;
input 	loanio_gpio_loanio1_o_24;
input 	loanio_gpio_loanio1_o_25;
input 	loanio_gpio_loanio1_o_26;
input 	loanio_gpio_loanio1_o_27;
input 	loanio_gpio_loanio1_o_28;
input 	loanio_gpio_loanio2_o_0;
input 	loanio_gpio_loanio2_o_1;
input 	loanio_gpio_loanio2_o_2;
input 	loanio_gpio_loanio2_o_3;
input 	loanio_gpio_loanio2_o_4;
input 	loanio_gpio_loanio2_o_5;
input 	loanio_gpio_loanio2_o_6;
input 	loanio_gpio_loanio2_o_7;
input 	loanio_gpio_loanio2_o_8;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim0_inst;
output 	spim0_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_38;
output 	intermediate_39;
output 	uart0_inst;
output 	gpio_inst;
output 	gpio_inst1;
output 	gpio_inst2;
output 	gpio_inst3;
output 	gpio_inst4;
output 	gpio_inst5;
output 	gpio_inst6;
output 	gpio_inst7;
output 	gpio_inst8;
output 	gpio_inst9;
output 	gpio_inst10;
output 	gpio_inst11;
output 	gpio_inst12;
output 	gpio_inst13;
output 	gpio_inst14;
output 	gpio_inst15;
output 	gpio_inst16;
output 	gpio_inst17;
output 	gpio_inst18;
output 	gpio_inst19;
output 	gpio_inst20;
output 	gpio_inst21;
output 	gpio_inst22;
output 	gpio_inst23;
output 	gpio_inst24;
output 	gpio_inst25;
output 	gpio_inst26;
output 	gpio_inst27;
output 	gpio_inst28;
output 	gpio_inst29;
output 	gpio_inst30;
output 	gpio_inst31;
output 	gpio_inst32;
output 	gpio_inst33;
output 	gpio_inst34;
output 	gpio_inst35;
output 	gpio_inst36;
output 	gpio_inst37;
output 	gpio_inst38;
output 	gpio_inst39;
output 	gpio_inst40;
output 	gpio_inst41;
output 	gpio_inst42;
output 	gpio_inst43;
output 	gpio_inst44;
output 	gpio_inst45;
output 	gpio_inst46;
output 	gpio_inst47;
output 	gpio_inst48;
output 	gpio_inst49;
output 	gpio_inst50;
output 	gpio_inst51;
output 	gpio_inst52;
output 	gpio_inst53;
output 	gpio_inst54;
output 	gpio_inst55;
output 	gpio_inst56;
output 	gpio_inst57;
output 	gpio_inst58;
output 	gpio_inst59;
output 	gpio_inst60;
output 	gpio_inst61;
output 	gpio_inst62;
output 	gpio_inst63;
output 	gpio_inst64;
output 	gpio_inst65;
output 	gpio_inst66;
output 	intermediate_50;
output 	intermediate_40;
output 	intermediate_51;
output 	intermediate_41;
output 	intermediate_42;
output 	intermediate_52;
output 	intermediate_44;
output 	intermediate_54;
output 	intermediate_56;
output 	intermediate_58;
output 	intermediate_60;
output 	intermediate_62;
output 	intermediate_64;
output 	intermediate_43;
output 	intermediate_53;
output 	intermediate_45;
output 	intermediate_55;
output 	intermediate_57;
output 	intermediate_59;
output 	intermediate_61;
output 	intermediate_63;
output 	intermediate_65;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_47;
output 	intermediate_49;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_gpio_inst_GPIO62_0;
input 	hps_io_gpio_inst_LOANIO00_0;
input 	hps_io_gpio_inst_LOANIO41_0;
input 	hps_io_gpio_inst_LOANIO51_0;
input 	hps_io_gpio_inst_LOANIO52_0;
input 	hps_io_gpio_inst_LOANIO53_0;
input 	hps_io_gpio_inst_LOANIO54_0;
input 	hps_io_gpio_inst_LOANIO55_0;
input 	hps_io_gpio_inst_LOANIO56_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim0_inst_MISO;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_soc_system_hps_0_hps_io_border border(
	.gpio_loanio_loanio0_oe({loanio_gpio_loanio0_oe_28,loanio_gpio_loanio0_oe_27,loanio_gpio_loanio0_oe_26,loanio_gpio_loanio0_oe_25,loanio_gpio_loanio0_oe_24,loanio_gpio_loanio0_oe_23,loanio_gpio_loanio0_oe_22,loanio_gpio_loanio0_oe_21,loanio_gpio_loanio0_oe_20,loanio_gpio_loanio0_oe_19,
loanio_gpio_loanio0_oe_18,loanio_gpio_loanio0_oe_17,loanio_gpio_loanio0_oe_16,loanio_gpio_loanio0_oe_15,loanio_gpio_loanio0_oe_14,loanio_gpio_loanio0_oe_13,loanio_gpio_loanio0_oe_12,loanio_gpio_loanio0_oe_11,loanio_gpio_loanio0_oe_10,loanio_gpio_loanio0_oe_9,
loanio_gpio_loanio0_oe_8,loanio_gpio_loanio0_oe_7,loanio_gpio_loanio0_oe_6,loanio_gpio_loanio0_oe_5,loanio_gpio_loanio0_oe_4,loanio_gpio_loanio0_oe_3,loanio_gpio_loanio0_oe_2,loanio_gpio_loanio0_oe_1,loanio_gpio_loanio0_oe_0}),
	.gpio_loanio_loanio1_oe({loanio_gpio_loanio1_oe_28,loanio_gpio_loanio1_oe_27,loanio_gpio_loanio1_oe_26,loanio_gpio_loanio1_oe_25,loanio_gpio_loanio1_oe_24,loanio_gpio_loanio1_oe_23,loanio_gpio_loanio1_oe_22,loanio_gpio_loanio1_oe_21,loanio_gpio_loanio1_oe_20,loanio_gpio_loanio1_oe_19,
loanio_gpio_loanio1_oe_18,loanio_gpio_loanio1_oe_17,loanio_gpio_loanio1_oe_16,loanio_gpio_loanio1_oe_15,loanio_gpio_loanio1_oe_14,loanio_gpio_loanio1_oe_13,loanio_gpio_loanio1_oe_12,loanio_gpio_loanio1_oe_11,loanio_gpio_loanio1_oe_10,loanio_gpio_loanio1_oe_9,
loanio_gpio_loanio1_oe_8,loanio_gpio_loanio1_oe_7,loanio_gpio_loanio1_oe_6,loanio_gpio_loanio1_oe_5,loanio_gpio_loanio1_oe_4,loanio_gpio_loanio1_oe_3,loanio_gpio_loanio1_oe_2,loanio_gpio_loanio1_oe_1,loanio_gpio_loanio1_oe_0}),
	.gpio_loanio_loanio2_oe({loanio_gpio_loanio2_oe_8,loanio_gpio_loanio2_oe_7,loanio_gpio_loanio2_oe_6,loanio_gpio_loanio2_oe_5,loanio_gpio_loanio2_oe_4,loanio_gpio_loanio2_oe_3,loanio_gpio_loanio2_oe_2,loanio_gpio_loanio2_oe_1,loanio_gpio_loanio2_oe_0}),
	.gpio_loanio_loanio0_o({loanio_gpio_loanio0_o_28,loanio_gpio_loanio0_o_27,loanio_gpio_loanio0_o_26,loanio_gpio_loanio0_o_25,loanio_gpio_loanio0_o_24,loanio_gpio_loanio0_o_23,loanio_gpio_loanio0_o_22,loanio_gpio_loanio0_o_21,loanio_gpio_loanio0_o_20,loanio_gpio_loanio0_o_19,
loanio_gpio_loanio0_o_18,loanio_gpio_loanio0_o_17,loanio_gpio_loanio0_o_16,loanio_gpio_loanio0_o_15,loanio_gpio_loanio0_o_14,loanio_gpio_loanio0_o_13,loanio_gpio_loanio0_o_12,loanio_gpio_loanio0_o_11,loanio_gpio_loanio0_o_10,loanio_gpio_loanio0_o_9,
loanio_gpio_loanio0_o_8,loanio_gpio_loanio0_o_7,loanio_gpio_loanio0_o_6,loanio_gpio_loanio0_o_5,loanio_gpio_loanio0_o_4,loanio_gpio_loanio0_o_3,loanio_gpio_loanio0_o_2,loanio_gpio_loanio0_o_1,loanio_gpio_loanio0_o_0}),
	.gpio_loanio_loanio1_o({loanio_gpio_loanio1_o_28,loanio_gpio_loanio1_o_27,loanio_gpio_loanio1_o_26,loanio_gpio_loanio1_o_25,loanio_gpio_loanio1_o_24,loanio_gpio_loanio1_o_23,loanio_gpio_loanio1_o_22,loanio_gpio_loanio1_o_21,loanio_gpio_loanio1_o_20,loanio_gpio_loanio1_o_19,
loanio_gpio_loanio1_o_18,loanio_gpio_loanio1_o_17,loanio_gpio_loanio1_o_16,loanio_gpio_loanio1_o_15,loanio_gpio_loanio1_o_14,loanio_gpio_loanio1_o_13,loanio_gpio_loanio1_o_12,loanio_gpio_loanio1_o_11,loanio_gpio_loanio1_o_10,loanio_gpio_loanio1_o_9,
loanio_gpio_loanio1_o_8,loanio_gpio_loanio1_o_7,loanio_gpio_loanio1_o_6,loanio_gpio_loanio1_o_5,loanio_gpio_loanio1_o_4,loanio_gpio_loanio1_o_3,loanio_gpio_loanio1_o_2,loanio_gpio_loanio1_o_1,loanio_gpio_loanio1_o_0}),
	.gpio_loanio_loanio2_o({loanio_gpio_loanio2_o_8,loanio_gpio_loanio2_o_7,loanio_gpio_loanio2_o_6,loanio_gpio_loanio2_o_5,loanio_gpio_loanio2_o_4,loanio_gpio_loanio2_o_3,loanio_gpio_loanio2_o_2,loanio_gpio_loanio2_o_1,loanio_gpio_loanio2_o_0}),
	.hps_io_emac1_inst_TX_CLK({emac1_inst}),
	.hps_io_emac1_inst_TX_CTL({emac1_inst1}),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.hps_io_emac1_inst_MDC({emac1_inst2}),
	.hps_io_emac1_inst_TXD0({emac1_inst3}),
	.hps_io_emac1_inst_TXD1({emac1_inst4}),
	.hps_io_emac1_inst_TXD2({emac1_inst5}),
	.hps_io_emac1_inst_TXD3({emac1_inst6}),
	.hps_io_qspi_inst_CLK({qspi_inst}),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.hps_io_qspi_inst_SS0({qspi_inst1}),
	.hps_io_sdio_inst_CLK({sdio_inst}),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.hps_io_usb1_inst_STP({usb1_inst}),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.hps_io_spim0_inst_CLK({spim0_inst}),
	.hps_io_spim0_inst_SS0({spim0_inst1}),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.hps_io_spim1_inst_CLK({spim1_inst}),
	.hps_io_spim1_inst_SS0({spim1_inst1}),
	.intermediate_38(intermediate_38),
	.intermediate_39(intermediate_39),
	.hps_io_uart0_inst_TX({uart0_inst}),
	.gpio_loanio_loanio0_i({gpio_inst28,gpio_inst27,gpio_inst26,gpio_inst25,gpio_inst24,gpio_inst23,gpio_inst22,gpio_inst21,gpio_inst20,gpio_inst19,gpio_inst18,gpio_inst17,gpio_inst16,gpio_inst15,gpio_inst14,gpio_inst13,gpio_inst12,gpio_inst11,gpio_inst10,gpio_inst9,gpio_inst8,gpio_inst7,gpio_inst6,
gpio_inst5,gpio_inst4,gpio_inst3,gpio_inst2,gpio_inst1,gpio_inst}),
	.gpio_loanio_loanio1_i({gpio_inst57,gpio_inst56,gpio_inst55,gpio_inst54,gpio_inst53,gpio_inst52,gpio_inst51,gpio_inst50,gpio_inst49,gpio_inst48,gpio_inst47,gpio_inst46,gpio_inst45,gpio_inst44,gpio_inst43,gpio_inst42,gpio_inst41,gpio_inst40,gpio_inst39,gpio_inst38,gpio_inst37,gpio_inst36,gpio_inst35,
gpio_inst34,gpio_inst33,gpio_inst32,gpio_inst31,gpio_inst30,gpio_inst29}),
	.gpio_loanio_loanio2_i({gpio_inst66,gpio_inst65,gpio_inst64,gpio_inst63,gpio_inst62,gpio_inst61,gpio_inst60,gpio_inst59,gpio_inst58}),
	.intermediate_50(intermediate_50),
	.intermediate_40(intermediate_40),
	.intermediate_51(intermediate_51),
	.intermediate_41(intermediate_41),
	.intermediate_42(intermediate_42),
	.intermediate_52(intermediate_52),
	.intermediate_44(intermediate_44),
	.intermediate_54(intermediate_54),
	.intermediate_56(intermediate_56),
	.intermediate_58(intermediate_58),
	.intermediate_60(intermediate_60),
	.intermediate_62(intermediate_62),
	.intermediate_64(intermediate_64),
	.intermediate_43(intermediate_43),
	.intermediate_53(intermediate_53),
	.intermediate_45(intermediate_45),
	.intermediate_55(intermediate_55),
	.intermediate_57(intermediate_57),
	.intermediate_59(intermediate_59),
	.intermediate_61(intermediate_61),
	.intermediate_63(intermediate_63),
	.intermediate_65(intermediate_65),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_gpio_inst_GPIO62_0(hps_io_gpio_inst_GPIO62_0),
	.hps_io_gpio_inst_LOANIO00_0(hps_io_gpio_inst_LOANIO00_0),
	.hps_io_gpio_inst_LOANIO41_0(hps_io_gpio_inst_LOANIO41_0),
	.hps_io_gpio_inst_LOANIO51_0(hps_io_gpio_inst_LOANIO51_0),
	.hps_io_gpio_inst_LOANIO52_0(hps_io_gpio_inst_LOANIO52_0),
	.hps_io_gpio_inst_LOANIO53_0(hps_io_gpio_inst_LOANIO53_0),
	.hps_io_gpio_inst_LOANIO54_0(hps_io_gpio_inst_LOANIO54_0),
	.hps_io_gpio_inst_LOANIO55_0(hps_io_gpio_inst_LOANIO55_0),
	.hps_io_gpio_inst_LOANIO56_0(hps_io_gpio_inst_LOANIO56_0),
	.hps_io_emac1_inst_RXD0({hps_io_hps_io_emac1_inst_RXD0}),
	.hps_io_emac1_inst_RXD1({hps_io_hps_io_emac1_inst_RXD1}),
	.hps_io_emac1_inst_RXD2({hps_io_hps_io_emac1_inst_RXD2}),
	.hps_io_emac1_inst_RXD3({hps_io_hps_io_emac1_inst_RXD3}),
	.hps_io_emac1_inst_RX_CLK({hps_io_hps_io_emac1_inst_RX_CLK}),
	.hps_io_emac1_inst_RX_CTL({hps_io_hps_io_emac1_inst_RX_CTL}),
	.hps_io_spim0_inst_MISO({hps_io_hps_io_spim0_inst_MISO}),
	.hps_io_spim1_inst_MISO({hps_io_hps_io_spim1_inst_MISO}),
	.hps_io_uart0_inst_RX({hps_io_hps_io_uart0_inst_RX}),
	.hps_io_usb1_inst_CLK({hps_io_hps_io_usb1_inst_CLK}),
	.hps_io_usb1_inst_DIR({hps_io_hps_io_usb1_inst_DIR}),
	.hps_io_usb1_inst_NXT({hps_io_hps_io_usb1_inst_NXT}),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module soc_system_soc_system_hps_0_hps_io_border (
	gpio_loanio_loanio0_oe,
	gpio_loanio_loanio1_oe,
	gpio_loanio_loanio2_oe,
	gpio_loanio_loanio0_o,
	gpio_loanio_loanio1_o,
	gpio_loanio_loanio2_o,
	hps_io_emac1_inst_TX_CLK,
	hps_io_emac1_inst_TX_CTL,
	intermediate_0,
	intermediate_1,
	hps_io_emac1_inst_MDC,
	hps_io_emac1_inst_TXD0,
	hps_io_emac1_inst_TXD1,
	hps_io_emac1_inst_TXD2,
	hps_io_emac1_inst_TXD3,
	hps_io_qspi_inst_CLK,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	hps_io_qspi_inst_SS0,
	hps_io_sdio_inst_CLK,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	hps_io_usb1_inst_STP,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	hps_io_spim0_inst_CLK,
	hps_io_spim0_inst_SS0,
	intermediate_36,
	intermediate_37,
	hps_io_spim1_inst_CLK,
	hps_io_spim1_inst_SS0,
	intermediate_38,
	intermediate_39,
	hps_io_uart0_inst_TX,
	gpio_loanio_loanio0_i,
	gpio_loanio_loanio1_i,
	gpio_loanio_loanio2_i,
	intermediate_50,
	intermediate_40,
	intermediate_51,
	intermediate_41,
	intermediate_42,
	intermediate_52,
	intermediate_44,
	intermediate_54,
	intermediate_56,
	intermediate_58,
	intermediate_60,
	intermediate_62,
	intermediate_64,
	intermediate_43,
	intermediate_53,
	intermediate_45,
	intermediate_55,
	intermediate_57,
	intermediate_59,
	intermediate_61,
	intermediate_63,
	intermediate_65,
	intermediate_46,
	intermediate_48,
	intermediate_47,
	intermediate_49,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_gpio_inst_GPIO62_0,
	hps_io_gpio_inst_LOANIO00_0,
	hps_io_gpio_inst_LOANIO41_0,
	hps_io_gpio_inst_LOANIO51_0,
	hps_io_gpio_inst_LOANIO52_0,
	hps_io_gpio_inst_LOANIO53_0,
	hps_io_gpio_inst_LOANIO54_0,
	hps_io_gpio_inst_LOANIO55_0,
	hps_io_gpio_inst_LOANIO56_0,
	hps_io_emac1_inst_RXD0,
	hps_io_emac1_inst_RXD1,
	hps_io_emac1_inst_RXD2,
	hps_io_emac1_inst_RXD3,
	hps_io_emac1_inst_RX_CLK,
	hps_io_emac1_inst_RX_CTL,
	hps_io_spim0_inst_MISO,
	hps_io_spim1_inst_MISO,
	hps_io_uart0_inst_RX,
	hps_io_usb1_inst_CLK,
	hps_io_usb1_inst_DIR,
	hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
input 	[28:0] gpio_loanio_loanio0_oe;
input 	[28:0] gpio_loanio_loanio1_oe;
input 	[8:0] gpio_loanio_loanio2_oe;
input 	[28:0] gpio_loanio_loanio0_o;
input 	[28:0] gpio_loanio_loanio1_o;
input 	[8:0] gpio_loanio_loanio2_o;
output 	[0:0] hps_io_emac1_inst_TX_CLK;
output 	[0:0] hps_io_emac1_inst_TX_CTL;
output 	intermediate_0;
output 	intermediate_1;
output 	[0:0] hps_io_emac1_inst_MDC;
output 	[0:0] hps_io_emac1_inst_TXD0;
output 	[0:0] hps_io_emac1_inst_TXD1;
output 	[0:0] hps_io_emac1_inst_TXD2;
output 	[0:0] hps_io_emac1_inst_TXD3;
output 	[0:0] hps_io_qspi_inst_CLK;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	[0:0] hps_io_qspi_inst_SS0;
output 	[0:0] hps_io_sdio_inst_CLK;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	[0:0] hps_io_usb1_inst_STP;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	[0:0] hps_io_spim0_inst_CLK;
output 	[0:0] hps_io_spim0_inst_SS0;
output 	intermediate_36;
output 	intermediate_37;
output 	[0:0] hps_io_spim1_inst_CLK;
output 	[0:0] hps_io_spim1_inst_SS0;
output 	intermediate_38;
output 	intermediate_39;
output 	[0:0] hps_io_uart0_inst_TX;
output 	[28:0] gpio_loanio_loanio0_i;
output 	[28:0] gpio_loanio_loanio1_i;
output 	[8:0] gpio_loanio_loanio2_i;
output 	intermediate_50;
output 	intermediate_40;
output 	intermediate_51;
output 	intermediate_41;
output 	intermediate_42;
output 	intermediate_52;
output 	intermediate_44;
output 	intermediate_54;
output 	intermediate_56;
output 	intermediate_58;
output 	intermediate_60;
output 	intermediate_62;
output 	intermediate_64;
output 	intermediate_43;
output 	intermediate_53;
output 	intermediate_45;
output 	intermediate_55;
output 	intermediate_57;
output 	intermediate_59;
output 	intermediate_61;
output 	intermediate_63;
output 	intermediate_65;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_47;
output 	intermediate_49;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_gpio_inst_GPIO62_0;
input 	hps_io_gpio_inst_LOANIO00_0;
input 	hps_io_gpio_inst_LOANIO41_0;
input 	hps_io_gpio_inst_LOANIO51_0;
input 	hps_io_gpio_inst_LOANIO52_0;
input 	hps_io_gpio_inst_LOANIO53_0;
input 	hps_io_gpio_inst_LOANIO54_0;
input 	hps_io_gpio_inst_LOANIO55_0;
input 	hps_io_gpio_inst_LOANIO56_0;
input 	[0:0] hps_io_emac1_inst_RXD0;
input 	[0:0] hps_io_emac1_inst_RXD1;
input 	[0:0] hps_io_emac1_inst_RXD2;
input 	[0:0] hps_io_emac1_inst_RXD3;
input 	[0:0] hps_io_emac1_inst_RX_CLK;
input 	[0:0] hps_io_emac1_inst_RX_CTL;
input 	[0:0] hps_io_spim0_inst_MISO;
input 	[0:0] hps_io_spim1_inst_MISO;
input 	[0:0] hps_io_uart0_inst_RX;
input 	[0:0] hps_io_usb1_inst_CLK;
input 	[0:0] hps_io_usb1_inst_DIR;
input 	[0:0] hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdio_inst~O_SDMMC_PWR_EN ;
wire \uart0_inst~UARTRTSN ;
wire \~GND~combout ;

wire [3:0] emac1_inst_EMAC_PHY_TXD_bus;
wire [3:0] qspi_inst_QSPI_SS_N_bus;
wire [3:0] qspi_inst_QSPI_MO_EN_N_bus;
wire [7:0] sdio_inst_SDMMC_DATA_OE_bus;
wire [7:0] sdio_inst_SDMMC_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_OE_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_O_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_OE_bus;
wire [28:0] gpio_inst_LOANIO0_I_bus;
wire [28:0] gpio_inst_LOANIO1_I_bus;
wire [26:0] gpio_inst_LOANIO2_I_bus;

assign hps_io_emac1_inst_TXD0[0] = emac1_inst_EMAC_PHY_TXD_bus[0];
assign hps_io_emac1_inst_TXD1[0] = emac1_inst_EMAC_PHY_TXD_bus[1];
assign hps_io_emac1_inst_TXD2[0] = emac1_inst_EMAC_PHY_TXD_bus[2];
assign hps_io_emac1_inst_TXD3[0] = emac1_inst_EMAC_PHY_TXD_bus[3];

assign hps_io_qspi_inst_SS0[0] = qspi_inst_QSPI_SS_N_bus[0];

assign intermediate_3 = qspi_inst_QSPI_MO_EN_N_bus[0];
assign intermediate_5 = qspi_inst_QSPI_MO_EN_N_bus[1];
assign intermediate_7 = qspi_inst_QSPI_MO_EN_N_bus[2];
assign intermediate_9 = qspi_inst_QSPI_MO_EN_N_bus[3];

assign intermediate_13 = sdio_inst_SDMMC_DATA_OE_bus[0];
assign intermediate_15 = sdio_inst_SDMMC_DATA_OE_bus[1];
assign intermediate_17 = sdio_inst_SDMMC_DATA_OE_bus[2];
assign intermediate_19 = sdio_inst_SDMMC_DATA_OE_bus[3];

assign intermediate_12 = sdio_inst_SDMMC_DATA_O_bus[0];
assign intermediate_14 = sdio_inst_SDMMC_DATA_O_bus[1];
assign intermediate_16 = sdio_inst_SDMMC_DATA_O_bus[2];
assign intermediate_18 = sdio_inst_SDMMC_DATA_O_bus[3];

assign intermediate_20 = usb1_inst_USB_ULPI_DATA_O_bus[0];
assign intermediate_22 = usb1_inst_USB_ULPI_DATA_O_bus[1];
assign intermediate_24 = usb1_inst_USB_ULPI_DATA_O_bus[2];
assign intermediate_26 = usb1_inst_USB_ULPI_DATA_O_bus[3];
assign intermediate_28 = usb1_inst_USB_ULPI_DATA_O_bus[4];
assign intermediate_30 = usb1_inst_USB_ULPI_DATA_O_bus[5];
assign intermediate_32 = usb1_inst_USB_ULPI_DATA_O_bus[6];
assign intermediate_34 = usb1_inst_USB_ULPI_DATA_O_bus[7];

assign intermediate_21 = usb1_inst_USB_ULPI_DATA_OE_bus[0];
assign intermediate_23 = usb1_inst_USB_ULPI_DATA_OE_bus[1];
assign intermediate_25 = usb1_inst_USB_ULPI_DATA_OE_bus[2];
assign intermediate_27 = usb1_inst_USB_ULPI_DATA_OE_bus[3];
assign intermediate_29 = usb1_inst_USB_ULPI_DATA_OE_bus[4];
assign intermediate_31 = usb1_inst_USB_ULPI_DATA_OE_bus[5];
assign intermediate_33 = usb1_inst_USB_ULPI_DATA_OE_bus[6];
assign intermediate_35 = usb1_inst_USB_ULPI_DATA_OE_bus[7];

assign intermediate_42 = gpio_inst_GPIO1_PORTA_O_bus[11];
assign intermediate_52 = gpio_inst_GPIO1_PORTA_O_bus[12];
assign intermediate_44 = gpio_inst_GPIO1_PORTA_O_bus[19];
assign intermediate_54 = gpio_inst_GPIO1_PORTA_O_bus[22];
assign intermediate_56 = gpio_inst_GPIO1_PORTA_O_bus[23];
assign intermediate_58 = gpio_inst_GPIO1_PORTA_O_bus[24];
assign intermediate_60 = gpio_inst_GPIO1_PORTA_O_bus[25];
assign intermediate_62 = gpio_inst_GPIO1_PORTA_O_bus[26];
assign intermediate_64 = gpio_inst_GPIO1_PORTA_O_bus[27];

assign intermediate_51 = gpio_inst_GPIO0_PORTA_OE_bus[0];
assign intermediate_41 = gpio_inst_GPIO0_PORTA_OE_bus[9];

assign intermediate_46 = gpio_inst_GPIO2_PORTA_O_bus[3];
assign intermediate_48 = gpio_inst_GPIO2_PORTA_O_bus[4];

assign intermediate_50 = gpio_inst_GPIO0_PORTA_O_bus[0];
assign intermediate_40 = gpio_inst_GPIO0_PORTA_O_bus[9];

assign intermediate_47 = gpio_inst_GPIO2_PORTA_OE_bus[3];
assign intermediate_49 = gpio_inst_GPIO2_PORTA_OE_bus[4];

assign intermediate_43 = gpio_inst_GPIO1_PORTA_OE_bus[11];
assign intermediate_53 = gpio_inst_GPIO1_PORTA_OE_bus[12];
assign intermediate_45 = gpio_inst_GPIO1_PORTA_OE_bus[19];
assign intermediate_55 = gpio_inst_GPIO1_PORTA_OE_bus[22];
assign intermediate_57 = gpio_inst_GPIO1_PORTA_OE_bus[23];
assign intermediate_59 = gpio_inst_GPIO1_PORTA_OE_bus[24];
assign intermediate_61 = gpio_inst_GPIO1_PORTA_OE_bus[25];
assign intermediate_63 = gpio_inst_GPIO1_PORTA_OE_bus[26];
assign intermediate_65 = gpio_inst_GPIO1_PORTA_OE_bus[27];

assign gpio_loanio_loanio0_i[0] = gpio_inst_LOANIO0_I_bus[0];
assign gpio_loanio_loanio0_i[1] = gpio_inst_LOANIO0_I_bus[1];
assign gpio_loanio_loanio0_i[2] = gpio_inst_LOANIO0_I_bus[2];
assign gpio_loanio_loanio0_i[3] = gpio_inst_LOANIO0_I_bus[3];
assign gpio_loanio_loanio0_i[4] = gpio_inst_LOANIO0_I_bus[4];
assign gpio_loanio_loanio0_i[5] = gpio_inst_LOANIO0_I_bus[5];
assign gpio_loanio_loanio0_i[6] = gpio_inst_LOANIO0_I_bus[6];
assign gpio_loanio_loanio0_i[7] = gpio_inst_LOANIO0_I_bus[7];
assign gpio_loanio_loanio0_i[8] = gpio_inst_LOANIO0_I_bus[8];
assign gpio_loanio_loanio0_i[9] = gpio_inst_LOANIO0_I_bus[9];
assign gpio_loanio_loanio0_i[10] = gpio_inst_LOANIO0_I_bus[10];
assign gpio_loanio_loanio0_i[11] = gpio_inst_LOANIO0_I_bus[11];
assign gpio_loanio_loanio0_i[12] = gpio_inst_LOANIO0_I_bus[12];
assign gpio_loanio_loanio0_i[13] = gpio_inst_LOANIO0_I_bus[13];
assign gpio_loanio_loanio0_i[14] = gpio_inst_LOANIO0_I_bus[14];
assign gpio_loanio_loanio0_i[15] = gpio_inst_LOANIO0_I_bus[15];
assign gpio_loanio_loanio0_i[16] = gpio_inst_LOANIO0_I_bus[16];
assign gpio_loanio_loanio0_i[17] = gpio_inst_LOANIO0_I_bus[17];
assign gpio_loanio_loanio0_i[18] = gpio_inst_LOANIO0_I_bus[18];
assign gpio_loanio_loanio0_i[19] = gpio_inst_LOANIO0_I_bus[19];
assign gpio_loanio_loanio0_i[20] = gpio_inst_LOANIO0_I_bus[20];
assign gpio_loanio_loanio0_i[21] = gpio_inst_LOANIO0_I_bus[21];
assign gpio_loanio_loanio0_i[22] = gpio_inst_LOANIO0_I_bus[22];
assign gpio_loanio_loanio0_i[23] = gpio_inst_LOANIO0_I_bus[23];
assign gpio_loanio_loanio0_i[24] = gpio_inst_LOANIO0_I_bus[24];
assign gpio_loanio_loanio0_i[25] = gpio_inst_LOANIO0_I_bus[25];
assign gpio_loanio_loanio0_i[26] = gpio_inst_LOANIO0_I_bus[26];
assign gpio_loanio_loanio0_i[27] = gpio_inst_LOANIO0_I_bus[27];
assign gpio_loanio_loanio0_i[28] = gpio_inst_LOANIO0_I_bus[28];

assign gpio_loanio_loanio1_i[0] = gpio_inst_LOANIO1_I_bus[0];
assign gpio_loanio_loanio1_i[1] = gpio_inst_LOANIO1_I_bus[1];
assign gpio_loanio_loanio1_i[2] = gpio_inst_LOANIO1_I_bus[2];
assign gpio_loanio_loanio1_i[3] = gpio_inst_LOANIO1_I_bus[3];
assign gpio_loanio_loanio1_i[4] = gpio_inst_LOANIO1_I_bus[4];
assign gpio_loanio_loanio1_i[5] = gpio_inst_LOANIO1_I_bus[5];
assign gpio_loanio_loanio1_i[6] = gpio_inst_LOANIO1_I_bus[6];
assign gpio_loanio_loanio1_i[7] = gpio_inst_LOANIO1_I_bus[7];
assign gpio_loanio_loanio1_i[8] = gpio_inst_LOANIO1_I_bus[8];
assign gpio_loanio_loanio1_i[9] = gpio_inst_LOANIO1_I_bus[9];
assign gpio_loanio_loanio1_i[10] = gpio_inst_LOANIO1_I_bus[10];
assign gpio_loanio_loanio1_i[11] = gpio_inst_LOANIO1_I_bus[11];
assign gpio_loanio_loanio1_i[12] = gpio_inst_LOANIO1_I_bus[12];
assign gpio_loanio_loanio1_i[13] = gpio_inst_LOANIO1_I_bus[13];
assign gpio_loanio_loanio1_i[14] = gpio_inst_LOANIO1_I_bus[14];
assign gpio_loanio_loanio1_i[15] = gpio_inst_LOANIO1_I_bus[15];
assign gpio_loanio_loanio1_i[16] = gpio_inst_LOANIO1_I_bus[16];
assign gpio_loanio_loanio1_i[17] = gpio_inst_LOANIO1_I_bus[17];
assign gpio_loanio_loanio1_i[18] = gpio_inst_LOANIO1_I_bus[18];
assign gpio_loanio_loanio1_i[19] = gpio_inst_LOANIO1_I_bus[19];
assign gpio_loanio_loanio1_i[20] = gpio_inst_LOANIO1_I_bus[20];
assign gpio_loanio_loanio1_i[21] = gpio_inst_LOANIO1_I_bus[21];
assign gpio_loanio_loanio1_i[22] = gpio_inst_LOANIO1_I_bus[22];
assign gpio_loanio_loanio1_i[23] = gpio_inst_LOANIO1_I_bus[23];
assign gpio_loanio_loanio1_i[24] = gpio_inst_LOANIO1_I_bus[24];
assign gpio_loanio_loanio1_i[25] = gpio_inst_LOANIO1_I_bus[25];
assign gpio_loanio_loanio1_i[26] = gpio_inst_LOANIO1_I_bus[26];
assign gpio_loanio_loanio1_i[27] = gpio_inst_LOANIO1_I_bus[27];
assign gpio_loanio_loanio1_i[28] = gpio_inst_LOANIO1_I_bus[28];

assign gpio_loanio_loanio2_i[0] = gpio_inst_LOANIO2_I_bus[0];
assign gpio_loanio_loanio2_i[1] = gpio_inst_LOANIO2_I_bus[1];
assign gpio_loanio_loanio2_i[2] = gpio_inst_LOANIO2_I_bus[2];
assign gpio_loanio_loanio2_i[3] = gpio_inst_LOANIO2_I_bus[3];
assign gpio_loanio_loanio2_i[4] = gpio_inst_LOANIO2_I_bus[4];
assign gpio_loanio_loanio2_i[5] = gpio_inst_LOANIO2_I_bus[5];
assign gpio_loanio_loanio2_i[6] = gpio_inst_LOANIO2_I_bus[6];
assign gpio_loanio_loanio2_i[7] = gpio_inst_LOANIO2_I_bus[7];
assign gpio_loanio_loanio2_i[8] = gpio_inst_LOANIO2_I_bus[8];

soc_system_hps_sdram hps_sdram_inst(
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.GND_port(\~GND~combout ),
	.memory_oct_rzqin(memory_oct_rzqin));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_hps_peripheral_emac emac1_inst(
	.emac_clk_rx(hps_io_emac1_inst_RX_CLK[0]),
	.emac_phy_rxdv(hps_io_emac1_inst_RX_CTL[0]),
	.emac_gmii_mdo_i(hps_io_emac1_inst_MDIO_0),
	.emac_phy_rxd({hps_io_emac1_inst_RXD3[0],hps_io_emac1_inst_RXD2[0],hps_io_emac1_inst_RXD1[0],hps_io_emac1_inst_RXD0[0]}),
	.emac_clk_tx(hps_io_emac1_inst_TX_CLK[0]),
	.emac_phy_tx_oe(hps_io_emac1_inst_TX_CTL[0]),
	.emac_gmii_mdo_o(intermediate_0),
	.emac_gmii_mdo_oe(intermediate_1),
	.emac_gmii_mdc(hps_io_emac1_inst_MDC[0]),
	.emac_phy_txd(emac1_inst_EMAC_PHY_TXD_bus));
defparam emac1_inst.dummy_param = 256;

cyclonev_hps_peripheral_qspi qspi_inst(
	.qspi_mi0(hps_io_qspi_inst_IO0_0),
	.qspi_mi1(hps_io_qspi_inst_IO1_0),
	.qspi_mi2(hps_io_qspi_inst_IO2_0),
	.qspi_mi3(hps_io_qspi_inst_IO3_0),
	.qspi_sclk(hps_io_qspi_inst_CLK[0]),
	.qspi_mo0(intermediate_2),
	.qspi_mo1(intermediate_4),
	.qspi_mo2(intermediate_6),
	.qspi_mo3(intermediate_8),
	.qspi_mo_en_n(qspi_inst_QSPI_MO_EN_N_bus),
	.qspi_ss_n(qspi_inst_QSPI_SS_N_bus));
defparam qspi_inst.dummy_param = 256;

cyclonev_hps_peripheral_sdmmc sdio_inst(
	.sdmmc_fb_clk(gnd),
	.sdmmc_cmd_i(hps_io_sdio_inst_CMD_0),
	.sdmmc_data_i({gnd,gnd,gnd,gnd,hps_io_sdio_inst_D3_0,hps_io_sdio_inst_D2_0,hps_io_sdio_inst_D1_0,hps_io_sdio_inst_D0_0}),
	.sdmmc_pwr_en(\sdio_inst~O_SDMMC_PWR_EN ),
	.sdmmc_cclk(hps_io_sdio_inst_CLK[0]),
	.sdmmc_cmd_o(intermediate_10),
	.sdmmc_cmd_oe(intermediate_11),
	.sdmmc_data_o(sdio_inst_SDMMC_DATA_O_bus),
	.sdmmc_data_oe(sdio_inst_SDMMC_DATA_OE_bus));
defparam sdio_inst.dummy_param = 256;

cyclonev_hps_peripheral_usb usb1_inst(
	.usb_ulpi_clk(hps_io_usb1_inst_CLK[0]),
	.usb_ulpi_dir(hps_io_usb1_inst_DIR[0]),
	.usb_ulpi_nxt(hps_io_usb1_inst_NXT[0]),
	.usb_ulpi_data_i({hps_io_usb1_inst_D7_0,hps_io_usb1_inst_D6_0,hps_io_usb1_inst_D5_0,hps_io_usb1_inst_D4_0,hps_io_usb1_inst_D3_0,hps_io_usb1_inst_D2_0,hps_io_usb1_inst_D1_0,hps_io_usb1_inst_D0_0}),
	.usb_ulpi_stp(hps_io_usb1_inst_STP[0]),
	.usb_ulpi_data_o(usb1_inst_USB_ULPI_DATA_O_bus),
	.usb_ulpi_data_oe(usb1_inst_USB_ULPI_DATA_OE_bus));
defparam usb1_inst.dummy_param = 256;

cyclonev_hps_peripheral_spi_master spim0_inst(
	.spi_master_rxd(hps_io_spim0_inst_MISO[0]),
	.spi_master_sclk(hps_io_spim0_inst_CLK[0]),
	.spi_master_ss_0_n(hps_io_spim0_inst_SS0[0]),
	.spi_master_ss_1_n(),
	.spi_master_txd(intermediate_36),
	.spi_master_ssi_oe_n(intermediate_37));
defparam spim0_inst.dummy_param = 256;

cyclonev_hps_peripheral_spi_master spim1_inst(
	.spi_master_rxd(hps_io_spim1_inst_MISO[0]),
	.spi_master_sclk(hps_io_spim1_inst_CLK[0]),
	.spi_master_ss_0_n(hps_io_spim1_inst_SS0[0]),
	.spi_master_ss_1_n(),
	.spi_master_txd(intermediate_38),
	.spi_master_ssi_oe_n(intermediate_39));
defparam spim1_inst.dummy_param = 256;

cyclonev_hps_peripheral_uart uart0_inst(
	.uart_cts_n(gnd),
	.uart_rxd(hps_io_uart0_inst_RX[0]),
	.uart_rts_n(\uart0_inst~UARTRTSN ),
	.uart_txd(hps_io_uart0_inst_TX[0]));
defparam uart0_inst.dummy_param = 256;

cyclonev_hps_peripheral_gpio gpio_inst(
	.gpio0_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO09_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_LOANIO00_0}),
	.gpio1_porta_i({gnd,hps_io_gpio_inst_LOANIO56_0,hps_io_gpio_inst_LOANIO55_0,hps_io_gpio_inst_LOANIO54_0,hps_io_gpio_inst_LOANIO53_0,hps_io_gpio_inst_LOANIO52_0,hps_io_gpio_inst_LOANIO51_0,gnd,gnd,hps_io_gpio_inst_GPIO48_0,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_LOANIO41_0,
hps_io_gpio_inst_GPIO40_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.gpio2_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO62_0,hps_io_gpio_inst_GPIO61_0,gnd,gnd,gnd}),
	.loanio0_o({gpio_loanio_loanio0_o[28],gpio_loanio_loanio0_o[27],gpio_loanio_loanio0_o[26],gpio_loanio_loanio0_o[25],gpio_loanio_loanio0_o[24],gpio_loanio_loanio0_o[23],gpio_loanio_loanio0_o[22],gpio_loanio_loanio0_o[21],gpio_loanio_loanio0_o[20],gpio_loanio_loanio0_o[19],gpio_loanio_loanio0_o[18],gpio_loanio_loanio0_o[17],
gpio_loanio_loanio0_o[16],gpio_loanio_loanio0_o[15],gpio_loanio_loanio0_o[14],gpio_loanio_loanio0_o[13],gpio_loanio_loanio0_o[12],gpio_loanio_loanio0_o[11],gpio_loanio_loanio0_o[10],gpio_loanio_loanio0_o[9],gpio_loanio_loanio0_o[8],gpio_loanio_loanio0_o[7],gpio_loanio_loanio0_o[6],gpio_loanio_loanio0_o[5],
gpio_loanio_loanio0_o[4],gpio_loanio_loanio0_o[3],gpio_loanio_loanio0_o[2],gpio_loanio_loanio0_o[1],gpio_loanio_loanio0_o[0]}),
	.loanio0_oe({gpio_loanio_loanio0_oe[28],gpio_loanio_loanio0_oe[27],gpio_loanio_loanio0_oe[26],gpio_loanio_loanio0_oe[25],gpio_loanio_loanio0_oe[24],gpio_loanio_loanio0_oe[23],gpio_loanio_loanio0_oe[22],gpio_loanio_loanio0_oe[21],gpio_loanio_loanio0_oe[20],gpio_loanio_loanio0_oe[19],gpio_loanio_loanio0_oe[18],
gpio_loanio_loanio0_oe[17],gpio_loanio_loanio0_oe[16],gpio_loanio_loanio0_oe[15],gpio_loanio_loanio0_oe[14],gpio_loanio_loanio0_oe[13],gpio_loanio_loanio0_oe[12],gpio_loanio_loanio0_oe[11],gpio_loanio_loanio0_oe[10],gpio_loanio_loanio0_oe[9],gpio_loanio_loanio0_oe[8],gpio_loanio_loanio0_oe[7],
gpio_loanio_loanio0_oe[6],gpio_loanio_loanio0_oe[5],gpio_loanio_loanio0_oe[4],gpio_loanio_loanio0_oe[3],gpio_loanio_loanio0_oe[2],gpio_loanio_loanio0_oe[1],gpio_loanio_loanio0_oe[0]}),
	.loanio1_o({gpio_loanio_loanio1_o[28],gpio_loanio_loanio1_o[27],gpio_loanio_loanio1_o[26],gpio_loanio_loanio1_o[25],gpio_loanio_loanio1_o[24],gpio_loanio_loanio1_o[23],gpio_loanio_loanio1_o[22],gpio_loanio_loanio1_o[21],gpio_loanio_loanio1_o[20],gpio_loanio_loanio1_o[19],gpio_loanio_loanio1_o[18],gpio_loanio_loanio1_o[17],
gpio_loanio_loanio1_o[16],gpio_loanio_loanio1_o[15],gpio_loanio_loanio1_o[14],gpio_loanio_loanio1_o[13],gpio_loanio_loanio1_o[12],gpio_loanio_loanio1_o[11],gpio_loanio_loanio1_o[10],gpio_loanio_loanio1_o[9],gpio_loanio_loanio1_o[8],gpio_loanio_loanio1_o[7],gpio_loanio_loanio1_o[6],gpio_loanio_loanio1_o[5],
gpio_loanio_loanio1_o[4],gpio_loanio_loanio1_o[3],gpio_loanio_loanio1_o[2],gpio_loanio_loanio1_o[1],gpio_loanio_loanio1_o[0]}),
	.loanio1_oe({gpio_loanio_loanio1_oe[28],gpio_loanio_loanio1_oe[27],gpio_loanio_loanio1_oe[26],gpio_loanio_loanio1_oe[25],gpio_loanio_loanio1_oe[24],gpio_loanio_loanio1_oe[23],gpio_loanio_loanio1_oe[22],gpio_loanio_loanio1_oe[21],gpio_loanio_loanio1_oe[20],gpio_loanio_loanio1_oe[19],gpio_loanio_loanio1_oe[18],
gpio_loanio_loanio1_oe[17],gpio_loanio_loanio1_oe[16],gpio_loanio_loanio1_oe[15],gpio_loanio_loanio1_oe[14],gpio_loanio_loanio1_oe[13],gpio_loanio_loanio1_oe[12],gpio_loanio_loanio1_oe[11],gpio_loanio_loanio1_oe[10],gpio_loanio_loanio1_oe[9],gpio_loanio_loanio1_oe[8],gpio_loanio_loanio1_oe[7],
gpio_loanio_loanio1_oe[6],gpio_loanio_loanio1_oe[5],gpio_loanio_loanio1_oe[4],gpio_loanio_loanio1_oe[3],gpio_loanio_loanio1_oe[2],gpio_loanio_loanio1_oe[1],gpio_loanio_loanio1_oe[0]}),
	.loanio2_o({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gpio_loanio_loanio2_o[8],gpio_loanio_loanio2_o[7],gpio_loanio_loanio2_o[6],gpio_loanio_loanio2_o[5],gpio_loanio_loanio2_o[4],gpio_loanio_loanio2_o[3],gpio_loanio_loanio2_o[2],gpio_loanio_loanio2_o[1],gpio_loanio_loanio2_o[0]}),
	.loanio2_oe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gpio_loanio_loanio2_oe[8],gpio_loanio_loanio2_oe[7],gpio_loanio_loanio2_oe[6],gpio_loanio_loanio2_oe[5],gpio_loanio_loanio2_oe[4],gpio_loanio_loanio2_oe[3],gpio_loanio_loanio2_oe[2],gpio_loanio_loanio2_oe[1],
gpio_loanio_loanio2_oe[0]}),
	.loanio0_i(gpio_inst_LOANIO0_I_bus),
	.loanio1_i(gpio_inst_LOANIO1_I_bus),
	.loanio2_i(gpio_inst_LOANIO2_I_bus),
	.gpio0_porta_o(gpio_inst_GPIO0_PORTA_O_bus),
	.gpio0_porta_oe(gpio_inst_GPIO0_PORTA_OE_bus),
	.gpio1_porta_o(gpio_inst_GPIO1_PORTA_O_bus),
	.gpio1_porta_oe(gpio_inst_GPIO1_PORTA_OE_bus),
	.gpio2_porta_o(gpio_inst_GPIO2_PORTA_O_bus),
	.gpio2_porta_oe(gpio_inst_GPIO2_PORTA_OE_bus));
defparam gpio_inst.dummy_param = 256;

endmodule

module soc_system_hps_sdram (
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	GND_port,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	GND_port;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|afi_clk ;
wire \pll|pll_write_clk ;
wire \p0|umemphy|afi_cal_fail ;
wire \p0|umemphy|afi_cal_success ;
wire \p0|umemphy|afi_rdata_valid[0] ;
wire \p0|umemphy|ctl_reset_n ;
wire \p0|umemphy|afi_rdata[0] ;
wire \p0|umemphy|afi_rdata[1] ;
wire \p0|umemphy|afi_rdata[2] ;
wire \p0|umemphy|afi_rdata[3] ;
wire \p0|umemphy|afi_rdata[4] ;
wire \p0|umemphy|afi_rdata[5] ;
wire \p0|umemphy|afi_rdata[6] ;
wire \p0|umemphy|afi_rdata[7] ;
wire \p0|umemphy|afi_rdata[8] ;
wire \p0|umemphy|afi_rdata[9] ;
wire \p0|umemphy|afi_rdata[10] ;
wire \p0|umemphy|afi_rdata[11] ;
wire \p0|umemphy|afi_rdata[12] ;
wire \p0|umemphy|afi_rdata[13] ;
wire \p0|umemphy|afi_rdata[14] ;
wire \p0|umemphy|afi_rdata[15] ;
wire \p0|umemphy|afi_rdata[16] ;
wire \p0|umemphy|afi_rdata[17] ;
wire \p0|umemphy|afi_rdata[18] ;
wire \p0|umemphy|afi_rdata[19] ;
wire \p0|umemphy|afi_rdata[20] ;
wire \p0|umemphy|afi_rdata[21] ;
wire \p0|umemphy|afi_rdata[22] ;
wire \p0|umemphy|afi_rdata[23] ;
wire \p0|umemphy|afi_rdata[24] ;
wire \p0|umemphy|afi_rdata[25] ;
wire \p0|umemphy|afi_rdata[26] ;
wire \p0|umemphy|afi_rdata[27] ;
wire \p0|umemphy|afi_rdata[28] ;
wire \p0|umemphy|afi_rdata[29] ;
wire \p0|umemphy|afi_rdata[30] ;
wire \p0|umemphy|afi_rdata[31] ;
wire \p0|umemphy|afi_rdata[32] ;
wire \p0|umemphy|afi_rdata[33] ;
wire \p0|umemphy|afi_rdata[34] ;
wire \p0|umemphy|afi_rdata[35] ;
wire \p0|umemphy|afi_rdata[36] ;
wire \p0|umemphy|afi_rdata[37] ;
wire \p0|umemphy|afi_rdata[38] ;
wire \p0|umemphy|afi_rdata[39] ;
wire \p0|umemphy|afi_rdata[40] ;
wire \p0|umemphy|afi_rdata[41] ;
wire \p0|umemphy|afi_rdata[42] ;
wire \p0|umemphy|afi_rdata[43] ;
wire \p0|umemphy|afi_rdata[44] ;
wire \p0|umemphy|afi_rdata[45] ;
wire \p0|umemphy|afi_rdata[46] ;
wire \p0|umemphy|afi_rdata[47] ;
wire \p0|umemphy|afi_rdata[48] ;
wire \p0|umemphy|afi_rdata[49] ;
wire \p0|umemphy|afi_rdata[50] ;
wire \p0|umemphy|afi_rdata[51] ;
wire \p0|umemphy|afi_rdata[52] ;
wire \p0|umemphy|afi_rdata[53] ;
wire \p0|umemphy|afi_rdata[54] ;
wire \p0|umemphy|afi_rdata[55] ;
wire \p0|umemphy|afi_rdata[56] ;
wire \p0|umemphy|afi_rdata[57] ;
wire \p0|umemphy|afi_rdata[58] ;
wire \p0|umemphy|afi_rdata[59] ;
wire \p0|umemphy|afi_rdata[60] ;
wire \p0|umemphy|afi_rdata[61] ;
wire \p0|umemphy|afi_rdata[62] ;
wire \p0|umemphy|afi_rdata[63] ;
wire \p0|umemphy|afi_rdata[64] ;
wire \p0|umemphy|afi_rdata[65] ;
wire \p0|umemphy|afi_rdata[66] ;
wire \p0|umemphy|afi_rdata[67] ;
wire \p0|umemphy|afi_rdata[68] ;
wire \p0|umemphy|afi_rdata[69] ;
wire \p0|umemphy|afi_rdata[70] ;
wire \p0|umemphy|afi_rdata[71] ;
wire \p0|umemphy|afi_rdata[72] ;
wire \p0|umemphy|afi_rdata[73] ;
wire \p0|umemphy|afi_rdata[74] ;
wire \p0|umemphy|afi_rdata[75] ;
wire \p0|umemphy|afi_rdata[76] ;
wire \p0|umemphy|afi_rdata[77] ;
wire \p0|umemphy|afi_rdata[78] ;
wire \p0|umemphy|afi_rdata[79] ;
wire \p0|umemphy|afi_wlat[0] ;
wire \p0|umemphy|afi_wlat[1] ;
wire \p0|umemphy|afi_wlat[2] ;
wire \p0|umemphy|afi_wlat[3] ;
wire \c0|afi_cas_n[0] ;
wire \c0|afi_ras_n[0] ;
wire \c0|afi_rst_n[0] ;
wire \c0|afi_we_n[0] ;
wire \c0|afi_addr[0] ;
wire \c0|afi_addr[1] ;
wire \c0|afi_addr[2] ;
wire \c0|afi_addr[3] ;
wire \c0|afi_addr[4] ;
wire \c0|afi_addr[5] ;
wire \c0|afi_addr[6] ;
wire \c0|afi_addr[7] ;
wire \c0|afi_addr[8] ;
wire \c0|afi_addr[9] ;
wire \c0|afi_addr[10] ;
wire \c0|afi_addr[11] ;
wire \c0|afi_addr[12] ;
wire \c0|afi_addr[13] ;
wire \c0|afi_addr[14] ;
wire \c0|afi_addr[15] ;
wire \c0|afi_addr[16] ;
wire \c0|afi_addr[17] ;
wire \c0|afi_addr[18] ;
wire \c0|afi_addr[19] ;
wire \c0|afi_ba[0] ;
wire \c0|afi_ba[1] ;
wire \c0|afi_ba[2] ;
wire \c0|afi_cke[0] ;
wire \c0|afi_cke[1] ;
wire \c0|afi_cs_n[0] ;
wire \c0|afi_cs_n[1] ;
wire \c0|afi_dm_int[0] ;
wire \c0|afi_dm_int[1] ;
wire \c0|afi_dm_int[2] ;
wire \c0|afi_dm_int[3] ;
wire \c0|afi_dm_int[4] ;
wire \c0|afi_dm_int[5] ;
wire \c0|afi_dm_int[6] ;
wire \c0|afi_dm_int[7] ;
wire \c0|afi_dm_int[8] ;
wire \c0|afi_dm_int[9] ;
wire \c0|afi_dqs_burst[0] ;
wire \c0|afi_dqs_burst[1] ;
wire \c0|afi_dqs_burst[2] ;
wire \c0|afi_dqs_burst[3] ;
wire \c0|afi_dqs_burst[4] ;
wire \c0|afi_odt[0] ;
wire \c0|afi_odt[1] ;
wire \c0|afi_rdata_en[0] ;
wire \c0|afi_rdata_en[1] ;
wire \c0|afi_rdata_en[2] ;
wire \c0|afi_rdata_en[3] ;
wire \c0|afi_rdata_en[4] ;
wire \c0|afi_rdata_en_full[0] ;
wire \c0|afi_rdata_en_full[1] ;
wire \c0|afi_rdata_en_full[2] ;
wire \c0|afi_rdata_en_full[3] ;
wire \c0|afi_rdata_en_full[4] ;
wire \c0|afi_wdata_int[0] ;
wire \c0|afi_wdata_int[1] ;
wire \c0|afi_wdata_int[2] ;
wire \c0|afi_wdata_int[3] ;
wire \c0|afi_wdata_int[4] ;
wire \c0|afi_wdata_int[5] ;
wire \c0|afi_wdata_int[6] ;
wire \c0|afi_wdata_int[7] ;
wire \c0|afi_wdata_int[8] ;
wire \c0|afi_wdata_int[9] ;
wire \c0|afi_wdata_int[10] ;
wire \c0|afi_wdata_int[11] ;
wire \c0|afi_wdata_int[12] ;
wire \c0|afi_wdata_int[13] ;
wire \c0|afi_wdata_int[14] ;
wire \c0|afi_wdata_int[15] ;
wire \c0|afi_wdata_int[16] ;
wire \c0|afi_wdata_int[17] ;
wire \c0|afi_wdata_int[18] ;
wire \c0|afi_wdata_int[19] ;
wire \c0|afi_wdata_int[20] ;
wire \c0|afi_wdata_int[21] ;
wire \c0|afi_wdata_int[22] ;
wire \c0|afi_wdata_int[23] ;
wire \c0|afi_wdata_int[24] ;
wire \c0|afi_wdata_int[25] ;
wire \c0|afi_wdata_int[26] ;
wire \c0|afi_wdata_int[27] ;
wire \c0|afi_wdata_int[28] ;
wire \c0|afi_wdata_int[29] ;
wire \c0|afi_wdata_int[30] ;
wire \c0|afi_wdata_int[31] ;
wire \c0|afi_wdata_int[32] ;
wire \c0|afi_wdata_int[33] ;
wire \c0|afi_wdata_int[34] ;
wire \c0|afi_wdata_int[35] ;
wire \c0|afi_wdata_int[36] ;
wire \c0|afi_wdata_int[37] ;
wire \c0|afi_wdata_int[38] ;
wire \c0|afi_wdata_int[39] ;
wire \c0|afi_wdata_int[40] ;
wire \c0|afi_wdata_int[41] ;
wire \c0|afi_wdata_int[42] ;
wire \c0|afi_wdata_int[43] ;
wire \c0|afi_wdata_int[44] ;
wire \c0|afi_wdata_int[45] ;
wire \c0|afi_wdata_int[46] ;
wire \c0|afi_wdata_int[47] ;
wire \c0|afi_wdata_int[48] ;
wire \c0|afi_wdata_int[49] ;
wire \c0|afi_wdata_int[50] ;
wire \c0|afi_wdata_int[51] ;
wire \c0|afi_wdata_int[52] ;
wire \c0|afi_wdata_int[53] ;
wire \c0|afi_wdata_int[54] ;
wire \c0|afi_wdata_int[55] ;
wire \c0|afi_wdata_int[56] ;
wire \c0|afi_wdata_int[57] ;
wire \c0|afi_wdata_int[58] ;
wire \c0|afi_wdata_int[59] ;
wire \c0|afi_wdata_int[60] ;
wire \c0|afi_wdata_int[61] ;
wire \c0|afi_wdata_int[62] ;
wire \c0|afi_wdata_int[63] ;
wire \c0|afi_wdata_int[64] ;
wire \c0|afi_wdata_int[65] ;
wire \c0|afi_wdata_int[66] ;
wire \c0|afi_wdata_int[67] ;
wire \c0|afi_wdata_int[68] ;
wire \c0|afi_wdata_int[69] ;
wire \c0|afi_wdata_int[70] ;
wire \c0|afi_wdata_int[71] ;
wire \c0|afi_wdata_int[72] ;
wire \c0|afi_wdata_int[73] ;
wire \c0|afi_wdata_int[74] ;
wire \c0|afi_wdata_int[75] ;
wire \c0|afi_wdata_int[76] ;
wire \c0|afi_wdata_int[77] ;
wire \c0|afi_wdata_int[78] ;
wire \c0|afi_wdata_int[79] ;
wire \c0|afi_wdata_valid[0] ;
wire \c0|afi_wdata_valid[1] ;
wire \c0|afi_wdata_valid[2] ;
wire \c0|afi_wdata_valid[3] ;
wire \c0|afi_wdata_valid[4] ;
wire \c0|cfg_addlat_wire[0] ;
wire \c0|cfg_addlat_wire[1] ;
wire \c0|cfg_addlat_wire[2] ;
wire \c0|cfg_addlat_wire[3] ;
wire \c0|cfg_addlat_wire[4] ;
wire \c0|cfg_bankaddrwidth_wire[0] ;
wire \c0|cfg_bankaddrwidth_wire[1] ;
wire \c0|cfg_bankaddrwidth_wire[2] ;
wire \c0|cfg_caswrlat_wire[0] ;
wire \c0|cfg_caswrlat_wire[1] ;
wire \c0|cfg_caswrlat_wire[2] ;
wire \c0|cfg_caswrlat_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[0] ;
wire \c0|cfg_coladdrwidth_wire[1] ;
wire \c0|cfg_coladdrwidth_wire[2] ;
wire \c0|cfg_coladdrwidth_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[4] ;
wire \c0|cfg_csaddrwidth_wire[0] ;
wire \c0|cfg_csaddrwidth_wire[1] ;
wire \c0|cfg_csaddrwidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[0] ;
wire \c0|cfg_devicewidth_wire[1] ;
wire \c0|cfg_devicewidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[0] ;
wire \c0|cfg_interfacewidth_wire[1] ;
wire \c0|cfg_interfacewidth_wire[2] ;
wire \c0|cfg_interfacewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[4] ;
wire \c0|cfg_interfacewidth_wire[5] ;
wire \c0|cfg_interfacewidth_wire[6] ;
wire \c0|cfg_interfacewidth_wire[7] ;
wire \c0|cfg_rowaddrwidth_wire[0] ;
wire \c0|cfg_rowaddrwidth_wire[1] ;
wire \c0|cfg_rowaddrwidth_wire[2] ;
wire \c0|cfg_rowaddrwidth_wire[3] ;
wire \c0|cfg_rowaddrwidth_wire[4] ;
wire \c0|cfg_tcl_wire[0] ;
wire \c0|cfg_tcl_wire[1] ;
wire \c0|cfg_tcl_wire[2] ;
wire \c0|cfg_tcl_wire[3] ;
wire \c0|cfg_tcl_wire[4] ;
wire \c0|cfg_tmrd_wire[0] ;
wire \c0|cfg_tmrd_wire[1] ;
wire \c0|cfg_tmrd_wire[2] ;
wire \c0|cfg_tmrd_wire[3] ;
wire \c0|cfg_trefi_wire[0] ;
wire \c0|cfg_trefi_wire[1] ;
wire \c0|cfg_trefi_wire[2] ;
wire \c0|cfg_trefi_wire[3] ;
wire \c0|cfg_trefi_wire[4] ;
wire \c0|cfg_trefi_wire[5] ;
wire \c0|cfg_trefi_wire[6] ;
wire \c0|cfg_trefi_wire[7] ;
wire \c0|cfg_trefi_wire[8] ;
wire \c0|cfg_trefi_wire[9] ;
wire \c0|cfg_trefi_wire[10] ;
wire \c0|cfg_trefi_wire[11] ;
wire \c0|cfg_trefi_wire[12] ;
wire \c0|cfg_trfc_wire[0] ;
wire \c0|cfg_trfc_wire[1] ;
wire \c0|cfg_trfc_wire[2] ;
wire \c0|cfg_trfc_wire[3] ;
wire \c0|cfg_trfc_wire[4] ;
wire \c0|cfg_trfc_wire[5] ;
wire \c0|cfg_trfc_wire[6] ;
wire \c0|cfg_trfc_wire[7] ;
wire \c0|cfg_twr_wire[0] ;
wire \c0|cfg_twr_wire[1] ;
wire \c0|cfg_twr_wire[2] ;
wire \c0|cfg_twr_wire[3] ;
wire \c0|afi_mem_clk_disable[0] ;
wire \c0|cfg_dramconfig_wire[0] ;
wire \c0|cfg_dramconfig_wire[1] ;
wire \c0|cfg_dramconfig_wire[2] ;
wire \c0|cfg_dramconfig_wire[3] ;
wire \c0|cfg_dramconfig_wire[4] ;
wire \c0|cfg_dramconfig_wire[5] ;
wire \c0|cfg_dramconfig_wire[6] ;
wire \c0|cfg_dramconfig_wire[7] ;
wire \c0|cfg_dramconfig_wire[8] ;
wire \c0|cfg_dramconfig_wire[9] ;
wire \c0|cfg_dramconfig_wire[10] ;
wire \c0|cfg_dramconfig_wire[11] ;
wire \c0|cfg_dramconfig_wire[12] ;
wire \c0|cfg_dramconfig_wire[13] ;
wire \c0|cfg_dramconfig_wire[14] ;
wire \c0|cfg_dramconfig_wire[15] ;
wire \c0|cfg_dramconfig_wire[16] ;
wire \c0|cfg_dramconfig_wire[17] ;
wire \c0|cfg_dramconfig_wire[18] ;
wire \c0|cfg_dramconfig_wire[19] ;
wire \c0|cfg_dramconfig_wire[20] ;
wire \p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ;
wire \dll|dll_delayctrl[0] ;
wire \dll|dll_delayctrl[1] ;
wire \dll|dll_delayctrl[2] ;
wire \dll|dll_delayctrl[3] ;
wire \dll|dll_delayctrl[4] ;
wire \dll|dll_delayctrl[5] ;
wire \dll|dll_delayctrl[6] ;


soc_system_hps_sdram_p0 p0(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid_0(\p0|umemphy|afi_rdata_valid[0] ),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata_0(\p0|umemphy|afi_rdata[0] ),
	.afi_rdata_1(\p0|umemphy|afi_rdata[1] ),
	.afi_rdata_2(\p0|umemphy|afi_rdata[2] ),
	.afi_rdata_3(\p0|umemphy|afi_rdata[3] ),
	.afi_rdata_4(\p0|umemphy|afi_rdata[4] ),
	.afi_rdata_5(\p0|umemphy|afi_rdata[5] ),
	.afi_rdata_6(\p0|umemphy|afi_rdata[6] ),
	.afi_rdata_7(\p0|umemphy|afi_rdata[7] ),
	.afi_rdata_8(\p0|umemphy|afi_rdata[8] ),
	.afi_rdata_9(\p0|umemphy|afi_rdata[9] ),
	.afi_rdata_10(\p0|umemphy|afi_rdata[10] ),
	.afi_rdata_11(\p0|umemphy|afi_rdata[11] ),
	.afi_rdata_12(\p0|umemphy|afi_rdata[12] ),
	.afi_rdata_13(\p0|umemphy|afi_rdata[13] ),
	.afi_rdata_14(\p0|umemphy|afi_rdata[14] ),
	.afi_rdata_15(\p0|umemphy|afi_rdata[15] ),
	.afi_rdata_16(\p0|umemphy|afi_rdata[16] ),
	.afi_rdata_17(\p0|umemphy|afi_rdata[17] ),
	.afi_rdata_18(\p0|umemphy|afi_rdata[18] ),
	.afi_rdata_19(\p0|umemphy|afi_rdata[19] ),
	.afi_rdata_20(\p0|umemphy|afi_rdata[20] ),
	.afi_rdata_21(\p0|umemphy|afi_rdata[21] ),
	.afi_rdata_22(\p0|umemphy|afi_rdata[22] ),
	.afi_rdata_23(\p0|umemphy|afi_rdata[23] ),
	.afi_rdata_24(\p0|umemphy|afi_rdata[24] ),
	.afi_rdata_25(\p0|umemphy|afi_rdata[25] ),
	.afi_rdata_26(\p0|umemphy|afi_rdata[26] ),
	.afi_rdata_27(\p0|umemphy|afi_rdata[27] ),
	.afi_rdata_28(\p0|umemphy|afi_rdata[28] ),
	.afi_rdata_29(\p0|umemphy|afi_rdata[29] ),
	.afi_rdata_30(\p0|umemphy|afi_rdata[30] ),
	.afi_rdata_31(\p0|umemphy|afi_rdata[31] ),
	.afi_rdata_32(\p0|umemphy|afi_rdata[32] ),
	.afi_rdata_33(\p0|umemphy|afi_rdata[33] ),
	.afi_rdata_34(\p0|umemphy|afi_rdata[34] ),
	.afi_rdata_35(\p0|umemphy|afi_rdata[35] ),
	.afi_rdata_36(\p0|umemphy|afi_rdata[36] ),
	.afi_rdata_37(\p0|umemphy|afi_rdata[37] ),
	.afi_rdata_38(\p0|umemphy|afi_rdata[38] ),
	.afi_rdata_39(\p0|umemphy|afi_rdata[39] ),
	.afi_rdata_40(\p0|umemphy|afi_rdata[40] ),
	.afi_rdata_41(\p0|umemphy|afi_rdata[41] ),
	.afi_rdata_42(\p0|umemphy|afi_rdata[42] ),
	.afi_rdata_43(\p0|umemphy|afi_rdata[43] ),
	.afi_rdata_44(\p0|umemphy|afi_rdata[44] ),
	.afi_rdata_45(\p0|umemphy|afi_rdata[45] ),
	.afi_rdata_46(\p0|umemphy|afi_rdata[46] ),
	.afi_rdata_47(\p0|umemphy|afi_rdata[47] ),
	.afi_rdata_48(\p0|umemphy|afi_rdata[48] ),
	.afi_rdata_49(\p0|umemphy|afi_rdata[49] ),
	.afi_rdata_50(\p0|umemphy|afi_rdata[50] ),
	.afi_rdata_51(\p0|umemphy|afi_rdata[51] ),
	.afi_rdata_52(\p0|umemphy|afi_rdata[52] ),
	.afi_rdata_53(\p0|umemphy|afi_rdata[53] ),
	.afi_rdata_54(\p0|umemphy|afi_rdata[54] ),
	.afi_rdata_55(\p0|umemphy|afi_rdata[55] ),
	.afi_rdata_56(\p0|umemphy|afi_rdata[56] ),
	.afi_rdata_57(\p0|umemphy|afi_rdata[57] ),
	.afi_rdata_58(\p0|umemphy|afi_rdata[58] ),
	.afi_rdata_59(\p0|umemphy|afi_rdata[59] ),
	.afi_rdata_60(\p0|umemphy|afi_rdata[60] ),
	.afi_rdata_61(\p0|umemphy|afi_rdata[61] ),
	.afi_rdata_62(\p0|umemphy|afi_rdata[62] ),
	.afi_rdata_63(\p0|umemphy|afi_rdata[63] ),
	.afi_rdata_64(\p0|umemphy|afi_rdata[64] ),
	.afi_rdata_65(\p0|umemphy|afi_rdata[65] ),
	.afi_rdata_66(\p0|umemphy|afi_rdata[66] ),
	.afi_rdata_67(\p0|umemphy|afi_rdata[67] ),
	.afi_rdata_68(\p0|umemphy|afi_rdata[68] ),
	.afi_rdata_69(\p0|umemphy|afi_rdata[69] ),
	.afi_rdata_70(\p0|umemphy|afi_rdata[70] ),
	.afi_rdata_71(\p0|umemphy|afi_rdata[71] ),
	.afi_rdata_72(\p0|umemphy|afi_rdata[72] ),
	.afi_rdata_73(\p0|umemphy|afi_rdata[73] ),
	.afi_rdata_74(\p0|umemphy|afi_rdata[74] ),
	.afi_rdata_75(\p0|umemphy|afi_rdata[75] ),
	.afi_rdata_76(\p0|umemphy|afi_rdata[76] ),
	.afi_rdata_77(\p0|umemphy|afi_rdata[77] ),
	.afi_rdata_78(\p0|umemphy|afi_rdata[78] ),
	.afi_rdata_79(\p0|umemphy|afi_rdata[79] ),
	.afi_wlat_0(\p0|umemphy|afi_wlat[0] ),
	.afi_wlat_1(\p0|umemphy|afi_wlat[1] ),
	.afi_wlat_2(\p0|umemphy|afi_wlat[2] ),
	.afi_wlat_3(\p0|umemphy|afi_wlat[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n_0(\c0|afi_cas_n[0] ),
	.afi_ras_n_0(\c0|afi_ras_n[0] ),
	.afi_rst_n_0(\c0|afi_rst_n[0] ),
	.afi_we_n_0(\c0|afi_we_n[0] ),
	.afi_addr_0(\c0|afi_addr[0] ),
	.afi_addr_1(\c0|afi_addr[1] ),
	.afi_addr_2(\c0|afi_addr[2] ),
	.afi_addr_3(\c0|afi_addr[3] ),
	.afi_addr_4(\c0|afi_addr[4] ),
	.afi_addr_5(\c0|afi_addr[5] ),
	.afi_addr_6(\c0|afi_addr[6] ),
	.afi_addr_7(\c0|afi_addr[7] ),
	.afi_addr_8(\c0|afi_addr[8] ),
	.afi_addr_9(\c0|afi_addr[9] ),
	.afi_addr_10(\c0|afi_addr[10] ),
	.afi_addr_11(\c0|afi_addr[11] ),
	.afi_addr_12(\c0|afi_addr[12] ),
	.afi_addr_13(\c0|afi_addr[13] ),
	.afi_addr_14(\c0|afi_addr[14] ),
	.afi_addr_15(\c0|afi_addr[15] ),
	.afi_addr_16(\c0|afi_addr[16] ),
	.afi_addr_17(\c0|afi_addr[17] ),
	.afi_addr_18(\c0|afi_addr[18] ),
	.afi_addr_19(\c0|afi_addr[19] ),
	.afi_ba_0(\c0|afi_ba[0] ),
	.afi_ba_1(\c0|afi_ba[1] ),
	.afi_ba_2(\c0|afi_ba[2] ),
	.afi_cke_0(\c0|afi_cke[0] ),
	.afi_cke_1(\c0|afi_cke[1] ),
	.afi_cs_n_0(\c0|afi_cs_n[0] ),
	.afi_cs_n_1(\c0|afi_cs_n[1] ),
	.afi_dm_int_0(\c0|afi_dm_int[0] ),
	.afi_dm_int_1(\c0|afi_dm_int[1] ),
	.afi_dm_int_2(\c0|afi_dm_int[2] ),
	.afi_dm_int_3(\c0|afi_dm_int[3] ),
	.afi_dm_int_4(\c0|afi_dm_int[4] ),
	.afi_dm_int_5(\c0|afi_dm_int[5] ),
	.afi_dm_int_6(\c0|afi_dm_int[6] ),
	.afi_dm_int_7(\c0|afi_dm_int[7] ),
	.afi_dm_int_8(\c0|afi_dm_int[8] ),
	.afi_dm_int_9(\c0|afi_dm_int[9] ),
	.afi_dqs_burst_0(\c0|afi_dqs_burst[0] ),
	.afi_dqs_burst_1(\c0|afi_dqs_burst[1] ),
	.afi_dqs_burst_2(\c0|afi_dqs_burst[2] ),
	.afi_dqs_burst_3(\c0|afi_dqs_burst[3] ),
	.afi_dqs_burst_4(\c0|afi_dqs_burst[4] ),
	.afi_odt_0(\c0|afi_odt[0] ),
	.afi_odt_1(\c0|afi_odt[1] ),
	.afi_rdata_en_0(\c0|afi_rdata_en[0] ),
	.afi_rdata_en_1(\c0|afi_rdata_en[1] ),
	.afi_rdata_en_2(\c0|afi_rdata_en[2] ),
	.afi_rdata_en_3(\c0|afi_rdata_en[3] ),
	.afi_rdata_en_4(\c0|afi_rdata_en[4] ),
	.afi_rdata_en_full_0(\c0|afi_rdata_en_full[0] ),
	.afi_rdata_en_full_1(\c0|afi_rdata_en_full[1] ),
	.afi_rdata_en_full_2(\c0|afi_rdata_en_full[2] ),
	.afi_rdata_en_full_3(\c0|afi_rdata_en_full[3] ),
	.afi_rdata_en_full_4(\c0|afi_rdata_en_full[4] ),
	.afi_wdata_int_0(\c0|afi_wdata_int[0] ),
	.afi_wdata_int_1(\c0|afi_wdata_int[1] ),
	.afi_wdata_int_2(\c0|afi_wdata_int[2] ),
	.afi_wdata_int_3(\c0|afi_wdata_int[3] ),
	.afi_wdata_int_4(\c0|afi_wdata_int[4] ),
	.afi_wdata_int_5(\c0|afi_wdata_int[5] ),
	.afi_wdata_int_6(\c0|afi_wdata_int[6] ),
	.afi_wdata_int_7(\c0|afi_wdata_int[7] ),
	.afi_wdata_int_8(\c0|afi_wdata_int[8] ),
	.afi_wdata_int_9(\c0|afi_wdata_int[9] ),
	.afi_wdata_int_10(\c0|afi_wdata_int[10] ),
	.afi_wdata_int_11(\c0|afi_wdata_int[11] ),
	.afi_wdata_int_12(\c0|afi_wdata_int[12] ),
	.afi_wdata_int_13(\c0|afi_wdata_int[13] ),
	.afi_wdata_int_14(\c0|afi_wdata_int[14] ),
	.afi_wdata_int_15(\c0|afi_wdata_int[15] ),
	.afi_wdata_int_16(\c0|afi_wdata_int[16] ),
	.afi_wdata_int_17(\c0|afi_wdata_int[17] ),
	.afi_wdata_int_18(\c0|afi_wdata_int[18] ),
	.afi_wdata_int_19(\c0|afi_wdata_int[19] ),
	.afi_wdata_int_20(\c0|afi_wdata_int[20] ),
	.afi_wdata_int_21(\c0|afi_wdata_int[21] ),
	.afi_wdata_int_22(\c0|afi_wdata_int[22] ),
	.afi_wdata_int_23(\c0|afi_wdata_int[23] ),
	.afi_wdata_int_24(\c0|afi_wdata_int[24] ),
	.afi_wdata_int_25(\c0|afi_wdata_int[25] ),
	.afi_wdata_int_26(\c0|afi_wdata_int[26] ),
	.afi_wdata_int_27(\c0|afi_wdata_int[27] ),
	.afi_wdata_int_28(\c0|afi_wdata_int[28] ),
	.afi_wdata_int_29(\c0|afi_wdata_int[29] ),
	.afi_wdata_int_30(\c0|afi_wdata_int[30] ),
	.afi_wdata_int_31(\c0|afi_wdata_int[31] ),
	.afi_wdata_int_32(\c0|afi_wdata_int[32] ),
	.afi_wdata_int_33(\c0|afi_wdata_int[33] ),
	.afi_wdata_int_34(\c0|afi_wdata_int[34] ),
	.afi_wdata_int_35(\c0|afi_wdata_int[35] ),
	.afi_wdata_int_36(\c0|afi_wdata_int[36] ),
	.afi_wdata_int_37(\c0|afi_wdata_int[37] ),
	.afi_wdata_int_38(\c0|afi_wdata_int[38] ),
	.afi_wdata_int_39(\c0|afi_wdata_int[39] ),
	.afi_wdata_int_40(\c0|afi_wdata_int[40] ),
	.afi_wdata_int_41(\c0|afi_wdata_int[41] ),
	.afi_wdata_int_42(\c0|afi_wdata_int[42] ),
	.afi_wdata_int_43(\c0|afi_wdata_int[43] ),
	.afi_wdata_int_44(\c0|afi_wdata_int[44] ),
	.afi_wdata_int_45(\c0|afi_wdata_int[45] ),
	.afi_wdata_int_46(\c0|afi_wdata_int[46] ),
	.afi_wdata_int_47(\c0|afi_wdata_int[47] ),
	.afi_wdata_int_48(\c0|afi_wdata_int[48] ),
	.afi_wdata_int_49(\c0|afi_wdata_int[49] ),
	.afi_wdata_int_50(\c0|afi_wdata_int[50] ),
	.afi_wdata_int_51(\c0|afi_wdata_int[51] ),
	.afi_wdata_int_52(\c0|afi_wdata_int[52] ),
	.afi_wdata_int_53(\c0|afi_wdata_int[53] ),
	.afi_wdata_int_54(\c0|afi_wdata_int[54] ),
	.afi_wdata_int_55(\c0|afi_wdata_int[55] ),
	.afi_wdata_int_56(\c0|afi_wdata_int[56] ),
	.afi_wdata_int_57(\c0|afi_wdata_int[57] ),
	.afi_wdata_int_58(\c0|afi_wdata_int[58] ),
	.afi_wdata_int_59(\c0|afi_wdata_int[59] ),
	.afi_wdata_int_60(\c0|afi_wdata_int[60] ),
	.afi_wdata_int_61(\c0|afi_wdata_int[61] ),
	.afi_wdata_int_62(\c0|afi_wdata_int[62] ),
	.afi_wdata_int_63(\c0|afi_wdata_int[63] ),
	.afi_wdata_int_64(\c0|afi_wdata_int[64] ),
	.afi_wdata_int_65(\c0|afi_wdata_int[65] ),
	.afi_wdata_int_66(\c0|afi_wdata_int[66] ),
	.afi_wdata_int_67(\c0|afi_wdata_int[67] ),
	.afi_wdata_int_68(\c0|afi_wdata_int[68] ),
	.afi_wdata_int_69(\c0|afi_wdata_int[69] ),
	.afi_wdata_int_70(\c0|afi_wdata_int[70] ),
	.afi_wdata_int_71(\c0|afi_wdata_int[71] ),
	.afi_wdata_int_72(\c0|afi_wdata_int[72] ),
	.afi_wdata_int_73(\c0|afi_wdata_int[73] ),
	.afi_wdata_int_74(\c0|afi_wdata_int[74] ),
	.afi_wdata_int_75(\c0|afi_wdata_int[75] ),
	.afi_wdata_int_76(\c0|afi_wdata_int[76] ),
	.afi_wdata_int_77(\c0|afi_wdata_int[77] ),
	.afi_wdata_int_78(\c0|afi_wdata_int[78] ),
	.afi_wdata_int_79(\c0|afi_wdata_int[79] ),
	.afi_wdata_valid_0(\c0|afi_wdata_valid[0] ),
	.afi_wdata_valid_1(\c0|afi_wdata_valid[1] ),
	.afi_wdata_valid_2(\c0|afi_wdata_valid[2] ),
	.afi_wdata_valid_3(\c0|afi_wdata_valid[3] ),
	.afi_wdata_valid_4(\c0|afi_wdata_valid[4] ),
	.cfg_addlat_wire_0(\c0|cfg_addlat_wire[0] ),
	.cfg_addlat_wire_1(\c0|cfg_addlat_wire[1] ),
	.cfg_addlat_wire_2(\c0|cfg_addlat_wire[2] ),
	.cfg_addlat_wire_3(\c0|cfg_addlat_wire[3] ),
	.cfg_addlat_wire_4(\c0|cfg_addlat_wire[4] ),
	.cfg_bankaddrwidth_wire_0(\c0|cfg_bankaddrwidth_wire[0] ),
	.cfg_bankaddrwidth_wire_1(\c0|cfg_bankaddrwidth_wire[1] ),
	.cfg_bankaddrwidth_wire_2(\c0|cfg_bankaddrwidth_wire[2] ),
	.cfg_caswrlat_wire_0(\c0|cfg_caswrlat_wire[0] ),
	.cfg_caswrlat_wire_1(\c0|cfg_caswrlat_wire[1] ),
	.cfg_caswrlat_wire_2(\c0|cfg_caswrlat_wire[2] ),
	.cfg_caswrlat_wire_3(\c0|cfg_caswrlat_wire[3] ),
	.cfg_coladdrwidth_wire_0(\c0|cfg_coladdrwidth_wire[0] ),
	.cfg_coladdrwidth_wire_1(\c0|cfg_coladdrwidth_wire[1] ),
	.cfg_coladdrwidth_wire_2(\c0|cfg_coladdrwidth_wire[2] ),
	.cfg_coladdrwidth_wire_3(\c0|cfg_coladdrwidth_wire[3] ),
	.cfg_coladdrwidth_wire_4(\c0|cfg_coladdrwidth_wire[4] ),
	.cfg_csaddrwidth_wire_0(\c0|cfg_csaddrwidth_wire[0] ),
	.cfg_csaddrwidth_wire_1(\c0|cfg_csaddrwidth_wire[1] ),
	.cfg_csaddrwidth_wire_2(\c0|cfg_csaddrwidth_wire[2] ),
	.cfg_devicewidth_wire_0(\c0|cfg_devicewidth_wire[0] ),
	.cfg_devicewidth_wire_1(\c0|cfg_devicewidth_wire[1] ),
	.cfg_devicewidth_wire_2(\c0|cfg_devicewidth_wire[2] ),
	.cfg_devicewidth_wire_3(\c0|cfg_devicewidth_wire[3] ),
	.cfg_interfacewidth_wire_0(\c0|cfg_interfacewidth_wire[0] ),
	.cfg_interfacewidth_wire_1(\c0|cfg_interfacewidth_wire[1] ),
	.cfg_interfacewidth_wire_2(\c0|cfg_interfacewidth_wire[2] ),
	.cfg_interfacewidth_wire_3(\c0|cfg_interfacewidth_wire[3] ),
	.cfg_interfacewidth_wire_4(\c0|cfg_interfacewidth_wire[4] ),
	.cfg_interfacewidth_wire_5(\c0|cfg_interfacewidth_wire[5] ),
	.cfg_interfacewidth_wire_6(\c0|cfg_interfacewidth_wire[6] ),
	.cfg_interfacewidth_wire_7(\c0|cfg_interfacewidth_wire[7] ),
	.cfg_rowaddrwidth_wire_0(\c0|cfg_rowaddrwidth_wire[0] ),
	.cfg_rowaddrwidth_wire_1(\c0|cfg_rowaddrwidth_wire[1] ),
	.cfg_rowaddrwidth_wire_2(\c0|cfg_rowaddrwidth_wire[2] ),
	.cfg_rowaddrwidth_wire_3(\c0|cfg_rowaddrwidth_wire[3] ),
	.cfg_rowaddrwidth_wire_4(\c0|cfg_rowaddrwidth_wire[4] ),
	.cfg_tcl_wire_0(\c0|cfg_tcl_wire[0] ),
	.cfg_tcl_wire_1(\c0|cfg_tcl_wire[1] ),
	.cfg_tcl_wire_2(\c0|cfg_tcl_wire[2] ),
	.cfg_tcl_wire_3(\c0|cfg_tcl_wire[3] ),
	.cfg_tcl_wire_4(\c0|cfg_tcl_wire[4] ),
	.cfg_tmrd_wire_0(\c0|cfg_tmrd_wire[0] ),
	.cfg_tmrd_wire_1(\c0|cfg_tmrd_wire[1] ),
	.cfg_tmrd_wire_2(\c0|cfg_tmrd_wire[2] ),
	.cfg_tmrd_wire_3(\c0|cfg_tmrd_wire[3] ),
	.cfg_trefi_wire_0(\c0|cfg_trefi_wire[0] ),
	.cfg_trefi_wire_1(\c0|cfg_trefi_wire[1] ),
	.cfg_trefi_wire_2(\c0|cfg_trefi_wire[2] ),
	.cfg_trefi_wire_3(\c0|cfg_trefi_wire[3] ),
	.cfg_trefi_wire_4(\c0|cfg_trefi_wire[4] ),
	.cfg_trefi_wire_5(\c0|cfg_trefi_wire[5] ),
	.cfg_trefi_wire_6(\c0|cfg_trefi_wire[6] ),
	.cfg_trefi_wire_7(\c0|cfg_trefi_wire[7] ),
	.cfg_trefi_wire_8(\c0|cfg_trefi_wire[8] ),
	.cfg_trefi_wire_9(\c0|cfg_trefi_wire[9] ),
	.cfg_trefi_wire_10(\c0|cfg_trefi_wire[10] ),
	.cfg_trefi_wire_11(\c0|cfg_trefi_wire[11] ),
	.cfg_trefi_wire_12(\c0|cfg_trefi_wire[12] ),
	.cfg_trfc_wire_0(\c0|cfg_trfc_wire[0] ),
	.cfg_trfc_wire_1(\c0|cfg_trfc_wire[1] ),
	.cfg_trfc_wire_2(\c0|cfg_trfc_wire[2] ),
	.cfg_trfc_wire_3(\c0|cfg_trfc_wire[3] ),
	.cfg_trfc_wire_4(\c0|cfg_trfc_wire[4] ),
	.cfg_trfc_wire_5(\c0|cfg_trfc_wire[5] ),
	.cfg_trfc_wire_6(\c0|cfg_trfc_wire[6] ),
	.cfg_trfc_wire_7(\c0|cfg_trfc_wire[7] ),
	.cfg_twr_wire_0(\c0|cfg_twr_wire[0] ),
	.cfg_twr_wire_1(\c0|cfg_twr_wire[1] ),
	.cfg_twr_wire_2(\c0|cfg_twr_wire[2] ),
	.cfg_twr_wire_3(\c0|cfg_twr_wire[3] ),
	.afi_mem_clk_disable_0(\c0|afi_mem_clk_disable[0] ),
	.cfg_dramconfig_wire_0(\c0|cfg_dramconfig_wire[0] ),
	.cfg_dramconfig_wire_1(\c0|cfg_dramconfig_wire[1] ),
	.cfg_dramconfig_wire_2(\c0|cfg_dramconfig_wire[2] ),
	.cfg_dramconfig_wire_3(\c0|cfg_dramconfig_wire[3] ),
	.cfg_dramconfig_wire_4(\c0|cfg_dramconfig_wire[4] ),
	.cfg_dramconfig_wire_5(\c0|cfg_dramconfig_wire[5] ),
	.cfg_dramconfig_wire_6(\c0|cfg_dramconfig_wire[6] ),
	.cfg_dramconfig_wire_7(\c0|cfg_dramconfig_wire[7] ),
	.cfg_dramconfig_wire_8(\c0|cfg_dramconfig_wire[8] ),
	.cfg_dramconfig_wire_9(\c0|cfg_dramconfig_wire[9] ),
	.cfg_dramconfig_wire_10(\c0|cfg_dramconfig_wire[10] ),
	.cfg_dramconfig_wire_11(\c0|cfg_dramconfig_wire[11] ),
	.cfg_dramconfig_wire_12(\c0|cfg_dramconfig_wire[12] ),
	.cfg_dramconfig_wire_13(\c0|cfg_dramconfig_wire[13] ),
	.cfg_dramconfig_wire_14(\c0|cfg_dramconfig_wire[14] ),
	.cfg_dramconfig_wire_15(\c0|cfg_dramconfig_wire[15] ),
	.cfg_dramconfig_wire_16(\c0|cfg_dramconfig_wire[16] ),
	.cfg_dramconfig_wire_17(\c0|cfg_dramconfig_wire[17] ),
	.cfg_dramconfig_wire_18(\c0|cfg_dramconfig_wire[18] ),
	.cfg_dramconfig_wire_19(\c0|cfg_dramconfig_wire[19] ),
	.cfg_dramconfig_wire_20(\c0|cfg_dramconfig_wire[20] ),
	.leveled_dqs_clocks_0(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ),
	.dll_delayctrl_0(\dll|dll_delayctrl[0] ),
	.dll_delayctrl_1(\dll|dll_delayctrl[1] ),
	.dll_delayctrl_2(\dll|dll_delayctrl[2] ),
	.dll_delayctrl_3(\dll|dll_delayctrl[3] ),
	.dll_delayctrl_4(\dll|dll_delayctrl[4] ),
	.dll_delayctrl_5(\dll|dll_delayctrl[5] ),
	.dll_delayctrl_6(\dll|dll_delayctrl[6] ),
	.GND_port(GND_port));

soc_system_hps_sdram_pll pll(
	.afi_half_clk(\pll|afi_clk ),
	.pll_write_clk_pre_phy_clk(\pll|pll_write_clk ));

soc_system_altera_mem_if_oct_cyclonev oct(
	.parallelterminationcontrol({parallelterminationcontrol_15,parallelterminationcontrol_14,parallelterminationcontrol_13,parallelterminationcontrol_12,parallelterminationcontrol_11,parallelterminationcontrol_10,parallelterminationcontrol_9,parallelterminationcontrol_8,
parallelterminationcontrol_7,parallelterminationcontrol_6,parallelterminationcontrol_5,parallelterminationcontrol_4,parallelterminationcontrol_3,parallelterminationcontrol_2,parallelterminationcontrol_1,parallelterminationcontrol_0}),
	.seriesterminationcontrol({seriesterminationcontrol_15,seriesterminationcontrol_14,seriesterminationcontrol_13,seriesterminationcontrol_12,seriesterminationcontrol_11,seriesterminationcontrol_10,seriesterminationcontrol_9,seriesterminationcontrol_8,seriesterminationcontrol_7,
seriesterminationcontrol_6,seriesterminationcontrol_5,seriesterminationcontrol_4,seriesterminationcontrol_3,seriesterminationcontrol_2,seriesterminationcontrol_1,seriesterminationcontrol_0}),
	.oct_rzqin(memory_oct_rzqin));

soc_system_altera_mem_if_dll_cyclonev dll(
	.clk(\pll|pll_write_clk ),
	.dll_delayctrl({\dll|dll_delayctrl[6] ,\dll|dll_delayctrl[5] ,\dll|dll_delayctrl[4] ,\dll|dll_delayctrl[3] ,\dll|dll_delayctrl[2] ,\dll|dll_delayctrl[1] ,\dll|dll_delayctrl[0] }));

soc_system_altera_mem_if_hard_memory_controller_top_cyclonev c0(
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid({\p0|umemphy|afi_rdata_valid[0] }),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata({\p0|umemphy|afi_rdata[79] ,\p0|umemphy|afi_rdata[78] ,\p0|umemphy|afi_rdata[77] ,\p0|umemphy|afi_rdata[76] ,\p0|umemphy|afi_rdata[75] ,\p0|umemphy|afi_rdata[74] ,\p0|umemphy|afi_rdata[73] ,\p0|umemphy|afi_rdata[72] ,\p0|umemphy|afi_rdata[71] ,
\p0|umemphy|afi_rdata[70] ,\p0|umemphy|afi_rdata[69] ,\p0|umemphy|afi_rdata[68] ,\p0|umemphy|afi_rdata[67] ,\p0|umemphy|afi_rdata[66] ,\p0|umemphy|afi_rdata[65] ,\p0|umemphy|afi_rdata[64] ,\p0|umemphy|afi_rdata[63] ,\p0|umemphy|afi_rdata[62] ,
\p0|umemphy|afi_rdata[61] ,\p0|umemphy|afi_rdata[60] ,\p0|umemphy|afi_rdata[59] ,\p0|umemphy|afi_rdata[58] ,\p0|umemphy|afi_rdata[57] ,\p0|umemphy|afi_rdata[56] ,\p0|umemphy|afi_rdata[55] ,\p0|umemphy|afi_rdata[54] ,\p0|umemphy|afi_rdata[53] ,
\p0|umemphy|afi_rdata[52] ,\p0|umemphy|afi_rdata[51] ,\p0|umemphy|afi_rdata[50] ,\p0|umemphy|afi_rdata[49] ,\p0|umemphy|afi_rdata[48] ,\p0|umemphy|afi_rdata[47] ,\p0|umemphy|afi_rdata[46] ,\p0|umemphy|afi_rdata[45] ,\p0|umemphy|afi_rdata[44] ,
\p0|umemphy|afi_rdata[43] ,\p0|umemphy|afi_rdata[42] ,\p0|umemphy|afi_rdata[41] ,\p0|umemphy|afi_rdata[40] ,\p0|umemphy|afi_rdata[39] ,\p0|umemphy|afi_rdata[38] ,\p0|umemphy|afi_rdata[37] ,\p0|umemphy|afi_rdata[36] ,\p0|umemphy|afi_rdata[35] ,
\p0|umemphy|afi_rdata[34] ,\p0|umemphy|afi_rdata[33] ,\p0|umemphy|afi_rdata[32] ,\p0|umemphy|afi_rdata[31] ,\p0|umemphy|afi_rdata[30] ,\p0|umemphy|afi_rdata[29] ,\p0|umemphy|afi_rdata[28] ,\p0|umemphy|afi_rdata[27] ,\p0|umemphy|afi_rdata[26] ,
\p0|umemphy|afi_rdata[25] ,\p0|umemphy|afi_rdata[24] ,\p0|umemphy|afi_rdata[23] ,\p0|umemphy|afi_rdata[22] ,\p0|umemphy|afi_rdata[21] ,\p0|umemphy|afi_rdata[20] ,\p0|umemphy|afi_rdata[19] ,\p0|umemphy|afi_rdata[18] ,\p0|umemphy|afi_rdata[17] ,
\p0|umemphy|afi_rdata[16] ,\p0|umemphy|afi_rdata[15] ,\p0|umemphy|afi_rdata[14] ,\p0|umemphy|afi_rdata[13] ,\p0|umemphy|afi_rdata[12] ,\p0|umemphy|afi_rdata[11] ,\p0|umemphy|afi_rdata[10] ,\p0|umemphy|afi_rdata[9] ,\p0|umemphy|afi_rdata[8] ,
\p0|umemphy|afi_rdata[7] ,\p0|umemphy|afi_rdata[6] ,\p0|umemphy|afi_rdata[5] ,\p0|umemphy|afi_rdata[4] ,\p0|umemphy|afi_rdata[3] ,\p0|umemphy|afi_rdata[2] ,\p0|umemphy|afi_rdata[1] ,\p0|umemphy|afi_rdata[0] }),
	.afi_wlat({\p0|umemphy|afi_wlat[3] ,\p0|umemphy|afi_wlat[2] ,\p0|umemphy|afi_wlat[1] ,\p0|umemphy|afi_wlat[0] }),
	.afi_cas_n({\c0|afi_cas_n[0] }),
	.afi_ras_n({\c0|afi_ras_n[0] }),
	.afi_rst_n({\c0|afi_rst_n[0] }),
	.afi_we_n({\c0|afi_we_n[0] }),
	.afi_addr({\c0|afi_addr[19] ,\c0|afi_addr[18] ,\c0|afi_addr[17] ,\c0|afi_addr[16] ,\c0|afi_addr[15] ,\c0|afi_addr[14] ,\c0|afi_addr[13] ,\c0|afi_addr[12] ,\c0|afi_addr[11] ,\c0|afi_addr[10] ,\c0|afi_addr[9] ,\c0|afi_addr[8] ,\c0|afi_addr[7] ,\c0|afi_addr[6] ,\c0|afi_addr[5] ,
\c0|afi_addr[4] ,\c0|afi_addr[3] ,\c0|afi_addr[2] ,\c0|afi_addr[1] ,\c0|afi_addr[0] }),
	.afi_ba({\c0|afi_ba[2] ,\c0|afi_ba[1] ,\c0|afi_ba[0] }),
	.afi_cke({\c0|afi_cke[1] ,\c0|afi_cke[0] }),
	.afi_cs_n({\c0|afi_cs_n[1] ,\c0|afi_cs_n[0] }),
	.afi_dm({\c0|afi_dm_int[9] ,\c0|afi_dm_int[8] ,\c0|afi_dm_int[7] ,\c0|afi_dm_int[6] ,\c0|afi_dm_int[5] ,\c0|afi_dm_int[4] ,\c0|afi_dm_int[3] ,\c0|afi_dm_int[2] ,\c0|afi_dm_int[1] ,\c0|afi_dm_int[0] }),
	.afi_dqs_burst({\c0|afi_dqs_burst[4] ,\c0|afi_dqs_burst[3] ,\c0|afi_dqs_burst[2] ,\c0|afi_dqs_burst[1] ,\c0|afi_dqs_burst[0] }),
	.afi_odt({\c0|afi_odt[1] ,\c0|afi_odt[0] }),
	.afi_rdata_en({\c0|afi_rdata_en[4] ,\c0|afi_rdata_en[3] ,\c0|afi_rdata_en[2] ,\c0|afi_rdata_en[1] ,\c0|afi_rdata_en[0] }),
	.afi_rdata_en_full({\c0|afi_rdata_en_full[4] ,\c0|afi_rdata_en_full[3] ,\c0|afi_rdata_en_full[2] ,\c0|afi_rdata_en_full[1] ,\c0|afi_rdata_en_full[0] }),
	.afi_wdata({\c0|afi_wdata_int[79] ,\c0|afi_wdata_int[78] ,\c0|afi_wdata_int[77] ,\c0|afi_wdata_int[76] ,\c0|afi_wdata_int[75] ,\c0|afi_wdata_int[74] ,\c0|afi_wdata_int[73] ,\c0|afi_wdata_int[72] ,\c0|afi_wdata_int[71] ,\c0|afi_wdata_int[70] ,\c0|afi_wdata_int[69] ,
\c0|afi_wdata_int[68] ,\c0|afi_wdata_int[67] ,\c0|afi_wdata_int[66] ,\c0|afi_wdata_int[65] ,\c0|afi_wdata_int[64] ,\c0|afi_wdata_int[63] ,\c0|afi_wdata_int[62] ,\c0|afi_wdata_int[61] ,\c0|afi_wdata_int[60] ,\c0|afi_wdata_int[59] ,\c0|afi_wdata_int[58] ,
\c0|afi_wdata_int[57] ,\c0|afi_wdata_int[56] ,\c0|afi_wdata_int[55] ,\c0|afi_wdata_int[54] ,\c0|afi_wdata_int[53] ,\c0|afi_wdata_int[52] ,\c0|afi_wdata_int[51] ,\c0|afi_wdata_int[50] ,\c0|afi_wdata_int[49] ,\c0|afi_wdata_int[48] ,\c0|afi_wdata_int[47] ,
\c0|afi_wdata_int[46] ,\c0|afi_wdata_int[45] ,\c0|afi_wdata_int[44] ,\c0|afi_wdata_int[43] ,\c0|afi_wdata_int[42] ,\c0|afi_wdata_int[41] ,\c0|afi_wdata_int[40] ,\c0|afi_wdata_int[39] ,\c0|afi_wdata_int[38] ,\c0|afi_wdata_int[37] ,\c0|afi_wdata_int[36] ,
\c0|afi_wdata_int[35] ,\c0|afi_wdata_int[34] ,\c0|afi_wdata_int[33] ,\c0|afi_wdata_int[32] ,\c0|afi_wdata_int[31] ,\c0|afi_wdata_int[30] ,\c0|afi_wdata_int[29] ,\c0|afi_wdata_int[28] ,\c0|afi_wdata_int[27] ,\c0|afi_wdata_int[26] ,\c0|afi_wdata_int[25] ,
\c0|afi_wdata_int[24] ,\c0|afi_wdata_int[23] ,\c0|afi_wdata_int[22] ,\c0|afi_wdata_int[21] ,\c0|afi_wdata_int[20] ,\c0|afi_wdata_int[19] ,\c0|afi_wdata_int[18] ,\c0|afi_wdata_int[17] ,\c0|afi_wdata_int[16] ,\c0|afi_wdata_int[15] ,\c0|afi_wdata_int[14] ,
\c0|afi_wdata_int[13] ,\c0|afi_wdata_int[12] ,\c0|afi_wdata_int[11] ,\c0|afi_wdata_int[10] ,\c0|afi_wdata_int[9] ,\c0|afi_wdata_int[8] ,\c0|afi_wdata_int[7] ,\c0|afi_wdata_int[6] ,\c0|afi_wdata_int[5] ,\c0|afi_wdata_int[4] ,\c0|afi_wdata_int[3] ,\c0|afi_wdata_int[2] ,
\c0|afi_wdata_int[1] ,\c0|afi_wdata_int[0] }),
	.afi_wdata_valid({\c0|afi_wdata_valid[4] ,\c0|afi_wdata_valid[3] ,\c0|afi_wdata_valid[2] ,\c0|afi_wdata_valid[1] ,\c0|afi_wdata_valid[0] }),
	.cfg_addlat({cfg_addlat_unconnected_wire_7,cfg_addlat_unconnected_wire_6,cfg_addlat_unconnected_wire_5,\c0|cfg_addlat_wire[4] ,\c0|cfg_addlat_wire[3] ,\c0|cfg_addlat_wire[2] ,\c0|cfg_addlat_wire[1] ,\c0|cfg_addlat_wire[0] }),
	.cfg_bankaddrwidth({cfg_bankaddrwidth_unconnected_wire_7,cfg_bankaddrwidth_unconnected_wire_6,cfg_bankaddrwidth_unconnected_wire_5,cfg_bankaddrwidth_unconnected_wire_4,cfg_bankaddrwidth_unconnected_wire_3,\c0|cfg_bankaddrwidth_wire[2] ,\c0|cfg_bankaddrwidth_wire[1] ,
\c0|cfg_bankaddrwidth_wire[0] }),
	.cfg_caswrlat({cfg_caswrlat_unconnected_wire_7,cfg_caswrlat_unconnected_wire_6,cfg_caswrlat_unconnected_wire_5,cfg_caswrlat_unconnected_wire_4,\c0|cfg_caswrlat_wire[3] ,\c0|cfg_caswrlat_wire[2] ,\c0|cfg_caswrlat_wire[1] ,\c0|cfg_caswrlat_wire[0] }),
	.cfg_coladdrwidth({cfg_coladdrwidth_unconnected_wire_7,cfg_coladdrwidth_unconnected_wire_6,cfg_coladdrwidth_unconnected_wire_5,\c0|cfg_coladdrwidth_wire[4] ,\c0|cfg_coladdrwidth_wire[3] ,\c0|cfg_coladdrwidth_wire[2] ,\c0|cfg_coladdrwidth_wire[1] ,\c0|cfg_coladdrwidth_wire[0] }),
	.cfg_csaddrwidth({cfg_csaddrwidth_unconnected_wire_7,cfg_csaddrwidth_unconnected_wire_6,cfg_csaddrwidth_unconnected_wire_5,cfg_csaddrwidth_unconnected_wire_4,cfg_csaddrwidth_unconnected_wire_3,\c0|cfg_csaddrwidth_wire[2] ,\c0|cfg_csaddrwidth_wire[1] ,\c0|cfg_csaddrwidth_wire[0] }),
	.cfg_devicewidth({cfg_devicewidth_unconnected_wire_7,cfg_devicewidth_unconnected_wire_6,cfg_devicewidth_unconnected_wire_5,cfg_devicewidth_unconnected_wire_4,\c0|cfg_devicewidth_wire[3] ,\c0|cfg_devicewidth_wire[2] ,\c0|cfg_devicewidth_wire[1] ,\c0|cfg_devicewidth_wire[0] }),
	.cfg_interfacewidth({\c0|cfg_interfacewidth_wire[7] ,\c0|cfg_interfacewidth_wire[6] ,\c0|cfg_interfacewidth_wire[5] ,\c0|cfg_interfacewidth_wire[4] ,\c0|cfg_interfacewidth_wire[3] ,\c0|cfg_interfacewidth_wire[2] ,\c0|cfg_interfacewidth_wire[1] ,\c0|cfg_interfacewidth_wire[0] }),
	.cfg_rowaddrwidth({cfg_rowaddrwidth_unconnected_wire_7,cfg_rowaddrwidth_unconnected_wire_6,cfg_rowaddrwidth_unconnected_wire_5,\c0|cfg_rowaddrwidth_wire[4] ,\c0|cfg_rowaddrwidth_wire[3] ,\c0|cfg_rowaddrwidth_wire[2] ,\c0|cfg_rowaddrwidth_wire[1] ,\c0|cfg_rowaddrwidth_wire[0] }),
	.cfg_tcl({cfg_tcl_unconnected_wire_7,cfg_tcl_unconnected_wire_6,cfg_tcl_unconnected_wire_5,\c0|cfg_tcl_wire[4] ,\c0|cfg_tcl_wire[3] ,\c0|cfg_tcl_wire[2] ,\c0|cfg_tcl_wire[1] ,\c0|cfg_tcl_wire[0] }),
	.cfg_tmrd({cfg_tmrd_unconnected_wire_7,cfg_tmrd_unconnected_wire_6,cfg_tmrd_unconnected_wire_5,cfg_tmrd_unconnected_wire_4,\c0|cfg_tmrd_wire[3] ,\c0|cfg_tmrd_wire[2] ,\c0|cfg_tmrd_wire[1] ,\c0|cfg_tmrd_wire[0] }),
	.cfg_trefi({cfg_trefi_unconnected_wire_15,cfg_trefi_unconnected_wire_14,cfg_trefi_unconnected_wire_13,\c0|cfg_trefi_wire[12] ,\c0|cfg_trefi_wire[11] ,\c0|cfg_trefi_wire[10] ,\c0|cfg_trefi_wire[9] ,\c0|cfg_trefi_wire[8] ,\c0|cfg_trefi_wire[7] ,\c0|cfg_trefi_wire[6] ,
\c0|cfg_trefi_wire[5] ,\c0|cfg_trefi_wire[4] ,\c0|cfg_trefi_wire[3] ,\c0|cfg_trefi_wire[2] ,\c0|cfg_trefi_wire[1] ,\c0|cfg_trefi_wire[0] }),
	.cfg_trfc({\c0|cfg_trfc_wire[7] ,\c0|cfg_trfc_wire[6] ,\c0|cfg_trfc_wire[5] ,\c0|cfg_trfc_wire[4] ,\c0|cfg_trfc_wire[3] ,\c0|cfg_trfc_wire[2] ,\c0|cfg_trfc_wire[1] ,\c0|cfg_trfc_wire[0] }),
	.cfg_twr({cfg_twr_unconnected_wire_7,cfg_twr_unconnected_wire_6,cfg_twr_unconnected_wire_5,cfg_twr_unconnected_wire_4,\c0|cfg_twr_wire[3] ,\c0|cfg_twr_wire[2] ,\c0|cfg_twr_wire[1] ,\c0|cfg_twr_wire[0] }),
	.afi_mem_clk_disable({\c0|afi_mem_clk_disable[0] }),
	.cfg_dramconfig({cfg_dramconfig_unconnected_wire_23,cfg_dramconfig_unconnected_wire_22,cfg_dramconfig_unconnected_wire_21,\c0|cfg_dramconfig_wire[20] ,\c0|cfg_dramconfig_wire[19] ,\c0|cfg_dramconfig_wire[18] ,\c0|cfg_dramconfig_wire[17] ,\c0|cfg_dramconfig_wire[16] ,
\c0|cfg_dramconfig_wire[15] ,\c0|cfg_dramconfig_wire[14] ,\c0|cfg_dramconfig_wire[13] ,\c0|cfg_dramconfig_wire[12] ,\c0|cfg_dramconfig_wire[11] ,\c0|cfg_dramconfig_wire[10] ,\c0|cfg_dramconfig_wire[9] ,\c0|cfg_dramconfig_wire[8] ,\c0|cfg_dramconfig_wire[7] ,
\c0|cfg_dramconfig_wire[6] ,\c0|cfg_dramconfig_wire[5] ,\c0|cfg_dramconfig_wire[4] ,\c0|cfg_dramconfig_wire[3] ,\c0|cfg_dramconfig_wire[2] ,\c0|cfg_dramconfig_wire[1] ,\c0|cfg_dramconfig_wire[0] }),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ));

endmodule

module soc_system_altera_mem_if_dll_cyclonev (
	clk,
	dll_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	[6:0] dll_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [6:0] dll_wys_m_DELAYCTRLOUT_bus;

assign dll_delayctrl[0] = dll_wys_m_DELAYCTRLOUT_bus[0];
assign dll_delayctrl[1] = dll_wys_m_DELAYCTRLOUT_bus[1];
assign dll_delayctrl[2] = dll_wys_m_DELAYCTRLOUT_bus[2];
assign dll_delayctrl[3] = dll_wys_m_DELAYCTRLOUT_bus[3];
assign dll_delayctrl[4] = dll_wys_m_DELAYCTRLOUT_bus[4];
assign dll_delayctrl[5] = dll_wys_m_DELAYCTRLOUT_bus[5];
assign dll_delayctrl[6] = dll_wys_m_DELAYCTRLOUT_bus[6];

cyclonev_dll dll_wys_m(
	.clk(clk),
	.aload(vcc),
	.upndnin(gnd),
	.upndninclkena(gnd),
	.dqsupdate(),
	.upndnout(),
	.delayctrlout(dll_wys_m_DELAYCTRLOUT_bus));
defparam dll_wys_m.delayctrlout_mode = "normal";
defparam dll_wys_m.input_frequency = "2500 ps";
defparam dll_wys_m.jitter_reduction = "true";
defparam dll_wys_m.sim_buffer_delay_increment = 10;
defparam dll_wys_m.sim_buffer_intrinsic_delay = 175;
defparam dll_wys_m.sim_valid_lock = 16;
defparam dll_wys_m.sim_valid_lockcount = 0;
defparam dll_wys_m.static_delay_ctrl = 8;
defparam dll_wys_m.upndnout_mode = "clock";
defparam dll_wys_m.use_upndnin = "false";
defparam dll_wys_m.use_upndninclkena = "false";

endmodule

module soc_system_altera_mem_if_hard_memory_controller_top_cyclonev (
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk)/* synthesis synthesis_greybox=0 */;
input 	afi_cal_fail;
input 	afi_cal_success;
input 	[0:0] afi_rdata_valid;
input 	ctl_reset_n;
input 	[79:0] afi_rdata;
input 	[3:0] afi_wlat;
output 	[0:0] afi_cas_n;
output 	[0:0] afi_ras_n;
output 	[0:0] afi_rst_n;
output 	[0:0] afi_we_n;
output 	[19:0] afi_addr;
output 	[2:0] afi_ba;
output 	[1:0] afi_cke;
output 	[1:0] afi_cs_n;
output 	[9:0] afi_dm;
output 	[4:0] afi_dqs_burst;
output 	[1:0] afi_odt;
output 	[4:0] afi_rdata_en;
output 	[4:0] afi_rdata_en_full;
output 	[79:0] afi_wdata;
output 	[4:0] afi_wdata_valid;
output 	[7:0] cfg_addlat;
output 	[7:0] cfg_bankaddrwidth;
output 	[7:0] cfg_caswrlat;
output 	[7:0] cfg_coladdrwidth;
output 	[7:0] cfg_csaddrwidth;
output 	[7:0] cfg_devicewidth;
output 	[7:0] cfg_interfacewidth;
output 	[7:0] cfg_rowaddrwidth;
output 	[7:0] cfg_tcl;
output 	[7:0] cfg_tmrd;
output 	[15:0] cfg_trefi;
output 	[7:0] cfg_trfc;
output 	[7:0] cfg_twr;
output 	[0:0] afi_mem_clk_disable;
output 	[23:0] cfg_dramconfig;
input 	ctl_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [19:0] hmc_inst_AFIADDR_bus;
wire [2:0] hmc_inst_AFIBA_bus;
wire [1:0] hmc_inst_AFICKE_bus;
wire [1:0] hmc_inst_AFICSN_bus;
wire [9:0] hmc_inst_AFIDM_bus;
wire [4:0] hmc_inst_AFIDQSBURST_bus;
wire [1:0] hmc_inst_AFIODT_bus;
wire [4:0] hmc_inst_AFIRDATAEN_bus;
wire [4:0] hmc_inst_AFIRDATAENFULL_bus;
wire [79:0] hmc_inst_AFIWDATA_bus;
wire [4:0] hmc_inst_AFIWDATAVALID_bus;
wire [4:0] hmc_inst_CFGADDLAT_bus;
wire [2:0] hmc_inst_CFGBANKADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGCASWRLAT_bus;
wire [4:0] hmc_inst_CFGCOLADDRWIDTH_bus;
wire [2:0] hmc_inst_CFGCSADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGDEVICEWIDTH_bus;
wire [7:0] hmc_inst_CFGINTERFACEWIDTH_bus;
wire [4:0] hmc_inst_CFGROWADDRWIDTH_bus;
wire [4:0] hmc_inst_CFGTCL_bus;
wire [3:0] hmc_inst_CFGTMRD_bus;
wire [12:0] hmc_inst_CFGTREFI_bus;
wire [7:0] hmc_inst_CFGTRFC_bus;
wire [3:0] hmc_inst_CFGTWR_bus;
wire [1:0] hmc_inst_CTLMEMCLKDISABLE_bus;
wire [20:0] hmc_inst_DRAMCONFIG_bus;

assign afi_addr[0] = hmc_inst_AFIADDR_bus[0];
assign afi_addr[1] = hmc_inst_AFIADDR_bus[1];
assign afi_addr[2] = hmc_inst_AFIADDR_bus[2];
assign afi_addr[3] = hmc_inst_AFIADDR_bus[3];
assign afi_addr[4] = hmc_inst_AFIADDR_bus[4];
assign afi_addr[5] = hmc_inst_AFIADDR_bus[5];
assign afi_addr[6] = hmc_inst_AFIADDR_bus[6];
assign afi_addr[7] = hmc_inst_AFIADDR_bus[7];
assign afi_addr[8] = hmc_inst_AFIADDR_bus[8];
assign afi_addr[9] = hmc_inst_AFIADDR_bus[9];
assign afi_addr[10] = hmc_inst_AFIADDR_bus[10];
assign afi_addr[11] = hmc_inst_AFIADDR_bus[11];
assign afi_addr[12] = hmc_inst_AFIADDR_bus[12];
assign afi_addr[13] = hmc_inst_AFIADDR_bus[13];
assign afi_addr[14] = hmc_inst_AFIADDR_bus[14];
assign afi_addr[15] = hmc_inst_AFIADDR_bus[15];
assign afi_addr[16] = hmc_inst_AFIADDR_bus[16];
assign afi_addr[17] = hmc_inst_AFIADDR_bus[17];
assign afi_addr[18] = hmc_inst_AFIADDR_bus[18];
assign afi_addr[19] = hmc_inst_AFIADDR_bus[19];

assign afi_ba[0] = hmc_inst_AFIBA_bus[0];
assign afi_ba[1] = hmc_inst_AFIBA_bus[1];
assign afi_ba[2] = hmc_inst_AFIBA_bus[2];

assign afi_cke[0] = hmc_inst_AFICKE_bus[0];
assign afi_cke[1] = hmc_inst_AFICKE_bus[1];

assign afi_cs_n[0] = hmc_inst_AFICSN_bus[0];
assign afi_cs_n[1] = hmc_inst_AFICSN_bus[1];

assign afi_dm[0] = hmc_inst_AFIDM_bus[0];
assign afi_dm[1] = hmc_inst_AFIDM_bus[1];
assign afi_dm[2] = hmc_inst_AFIDM_bus[2];
assign afi_dm[3] = hmc_inst_AFIDM_bus[3];
assign afi_dm[4] = hmc_inst_AFIDM_bus[4];
assign afi_dm[5] = hmc_inst_AFIDM_bus[5];
assign afi_dm[6] = hmc_inst_AFIDM_bus[6];
assign afi_dm[7] = hmc_inst_AFIDM_bus[7];
assign afi_dm[8] = hmc_inst_AFIDM_bus[8];
assign afi_dm[9] = hmc_inst_AFIDM_bus[9];

assign afi_dqs_burst[0] = hmc_inst_AFIDQSBURST_bus[0];
assign afi_dqs_burst[1] = hmc_inst_AFIDQSBURST_bus[1];
assign afi_dqs_burst[2] = hmc_inst_AFIDQSBURST_bus[2];
assign afi_dqs_burst[3] = hmc_inst_AFIDQSBURST_bus[3];
assign afi_dqs_burst[4] = hmc_inst_AFIDQSBURST_bus[4];

assign afi_odt[0] = hmc_inst_AFIODT_bus[0];
assign afi_odt[1] = hmc_inst_AFIODT_bus[1];

assign afi_rdata_en[0] = hmc_inst_AFIRDATAEN_bus[0];
assign afi_rdata_en[1] = hmc_inst_AFIRDATAEN_bus[1];
assign afi_rdata_en[2] = hmc_inst_AFIRDATAEN_bus[2];
assign afi_rdata_en[3] = hmc_inst_AFIRDATAEN_bus[3];
assign afi_rdata_en[4] = hmc_inst_AFIRDATAEN_bus[4];

assign afi_rdata_en_full[0] = hmc_inst_AFIRDATAENFULL_bus[0];
assign afi_rdata_en_full[1] = hmc_inst_AFIRDATAENFULL_bus[1];
assign afi_rdata_en_full[2] = hmc_inst_AFIRDATAENFULL_bus[2];
assign afi_rdata_en_full[3] = hmc_inst_AFIRDATAENFULL_bus[3];
assign afi_rdata_en_full[4] = hmc_inst_AFIRDATAENFULL_bus[4];

assign afi_wdata[0] = hmc_inst_AFIWDATA_bus[0];
assign afi_wdata[1] = hmc_inst_AFIWDATA_bus[1];
assign afi_wdata[2] = hmc_inst_AFIWDATA_bus[2];
assign afi_wdata[3] = hmc_inst_AFIWDATA_bus[3];
assign afi_wdata[4] = hmc_inst_AFIWDATA_bus[4];
assign afi_wdata[5] = hmc_inst_AFIWDATA_bus[5];
assign afi_wdata[6] = hmc_inst_AFIWDATA_bus[6];
assign afi_wdata[7] = hmc_inst_AFIWDATA_bus[7];
assign afi_wdata[8] = hmc_inst_AFIWDATA_bus[8];
assign afi_wdata[9] = hmc_inst_AFIWDATA_bus[9];
assign afi_wdata[10] = hmc_inst_AFIWDATA_bus[10];
assign afi_wdata[11] = hmc_inst_AFIWDATA_bus[11];
assign afi_wdata[12] = hmc_inst_AFIWDATA_bus[12];
assign afi_wdata[13] = hmc_inst_AFIWDATA_bus[13];
assign afi_wdata[14] = hmc_inst_AFIWDATA_bus[14];
assign afi_wdata[15] = hmc_inst_AFIWDATA_bus[15];
assign afi_wdata[16] = hmc_inst_AFIWDATA_bus[16];
assign afi_wdata[17] = hmc_inst_AFIWDATA_bus[17];
assign afi_wdata[18] = hmc_inst_AFIWDATA_bus[18];
assign afi_wdata[19] = hmc_inst_AFIWDATA_bus[19];
assign afi_wdata[20] = hmc_inst_AFIWDATA_bus[20];
assign afi_wdata[21] = hmc_inst_AFIWDATA_bus[21];
assign afi_wdata[22] = hmc_inst_AFIWDATA_bus[22];
assign afi_wdata[23] = hmc_inst_AFIWDATA_bus[23];
assign afi_wdata[24] = hmc_inst_AFIWDATA_bus[24];
assign afi_wdata[25] = hmc_inst_AFIWDATA_bus[25];
assign afi_wdata[26] = hmc_inst_AFIWDATA_bus[26];
assign afi_wdata[27] = hmc_inst_AFIWDATA_bus[27];
assign afi_wdata[28] = hmc_inst_AFIWDATA_bus[28];
assign afi_wdata[29] = hmc_inst_AFIWDATA_bus[29];
assign afi_wdata[30] = hmc_inst_AFIWDATA_bus[30];
assign afi_wdata[31] = hmc_inst_AFIWDATA_bus[31];
assign afi_wdata[32] = hmc_inst_AFIWDATA_bus[32];
assign afi_wdata[33] = hmc_inst_AFIWDATA_bus[33];
assign afi_wdata[34] = hmc_inst_AFIWDATA_bus[34];
assign afi_wdata[35] = hmc_inst_AFIWDATA_bus[35];
assign afi_wdata[36] = hmc_inst_AFIWDATA_bus[36];
assign afi_wdata[37] = hmc_inst_AFIWDATA_bus[37];
assign afi_wdata[38] = hmc_inst_AFIWDATA_bus[38];
assign afi_wdata[39] = hmc_inst_AFIWDATA_bus[39];
assign afi_wdata[40] = hmc_inst_AFIWDATA_bus[40];
assign afi_wdata[41] = hmc_inst_AFIWDATA_bus[41];
assign afi_wdata[42] = hmc_inst_AFIWDATA_bus[42];
assign afi_wdata[43] = hmc_inst_AFIWDATA_bus[43];
assign afi_wdata[44] = hmc_inst_AFIWDATA_bus[44];
assign afi_wdata[45] = hmc_inst_AFIWDATA_bus[45];
assign afi_wdata[46] = hmc_inst_AFIWDATA_bus[46];
assign afi_wdata[47] = hmc_inst_AFIWDATA_bus[47];
assign afi_wdata[48] = hmc_inst_AFIWDATA_bus[48];
assign afi_wdata[49] = hmc_inst_AFIWDATA_bus[49];
assign afi_wdata[50] = hmc_inst_AFIWDATA_bus[50];
assign afi_wdata[51] = hmc_inst_AFIWDATA_bus[51];
assign afi_wdata[52] = hmc_inst_AFIWDATA_bus[52];
assign afi_wdata[53] = hmc_inst_AFIWDATA_bus[53];
assign afi_wdata[54] = hmc_inst_AFIWDATA_bus[54];
assign afi_wdata[55] = hmc_inst_AFIWDATA_bus[55];
assign afi_wdata[56] = hmc_inst_AFIWDATA_bus[56];
assign afi_wdata[57] = hmc_inst_AFIWDATA_bus[57];
assign afi_wdata[58] = hmc_inst_AFIWDATA_bus[58];
assign afi_wdata[59] = hmc_inst_AFIWDATA_bus[59];
assign afi_wdata[60] = hmc_inst_AFIWDATA_bus[60];
assign afi_wdata[61] = hmc_inst_AFIWDATA_bus[61];
assign afi_wdata[62] = hmc_inst_AFIWDATA_bus[62];
assign afi_wdata[63] = hmc_inst_AFIWDATA_bus[63];
assign afi_wdata[64] = hmc_inst_AFIWDATA_bus[64];
assign afi_wdata[65] = hmc_inst_AFIWDATA_bus[65];
assign afi_wdata[66] = hmc_inst_AFIWDATA_bus[66];
assign afi_wdata[67] = hmc_inst_AFIWDATA_bus[67];
assign afi_wdata[68] = hmc_inst_AFIWDATA_bus[68];
assign afi_wdata[69] = hmc_inst_AFIWDATA_bus[69];
assign afi_wdata[70] = hmc_inst_AFIWDATA_bus[70];
assign afi_wdata[71] = hmc_inst_AFIWDATA_bus[71];
assign afi_wdata[72] = hmc_inst_AFIWDATA_bus[72];
assign afi_wdata[73] = hmc_inst_AFIWDATA_bus[73];
assign afi_wdata[74] = hmc_inst_AFIWDATA_bus[74];
assign afi_wdata[75] = hmc_inst_AFIWDATA_bus[75];
assign afi_wdata[76] = hmc_inst_AFIWDATA_bus[76];
assign afi_wdata[77] = hmc_inst_AFIWDATA_bus[77];
assign afi_wdata[78] = hmc_inst_AFIWDATA_bus[78];
assign afi_wdata[79] = hmc_inst_AFIWDATA_bus[79];

assign afi_wdata_valid[0] = hmc_inst_AFIWDATAVALID_bus[0];
assign afi_wdata_valid[1] = hmc_inst_AFIWDATAVALID_bus[1];
assign afi_wdata_valid[2] = hmc_inst_AFIWDATAVALID_bus[2];
assign afi_wdata_valid[3] = hmc_inst_AFIWDATAVALID_bus[3];
assign afi_wdata_valid[4] = hmc_inst_AFIWDATAVALID_bus[4];

assign cfg_addlat[0] = hmc_inst_CFGADDLAT_bus[0];
assign cfg_addlat[1] = hmc_inst_CFGADDLAT_bus[1];
assign cfg_addlat[2] = hmc_inst_CFGADDLAT_bus[2];
assign cfg_addlat[3] = hmc_inst_CFGADDLAT_bus[3];
assign cfg_addlat[4] = hmc_inst_CFGADDLAT_bus[4];

assign cfg_bankaddrwidth[0] = hmc_inst_CFGBANKADDRWIDTH_bus[0];
assign cfg_bankaddrwidth[1] = hmc_inst_CFGBANKADDRWIDTH_bus[1];
assign cfg_bankaddrwidth[2] = hmc_inst_CFGBANKADDRWIDTH_bus[2];

assign cfg_caswrlat[0] = hmc_inst_CFGCASWRLAT_bus[0];
assign cfg_caswrlat[1] = hmc_inst_CFGCASWRLAT_bus[1];
assign cfg_caswrlat[2] = hmc_inst_CFGCASWRLAT_bus[2];
assign cfg_caswrlat[3] = hmc_inst_CFGCASWRLAT_bus[3];

assign cfg_coladdrwidth[0] = hmc_inst_CFGCOLADDRWIDTH_bus[0];
assign cfg_coladdrwidth[1] = hmc_inst_CFGCOLADDRWIDTH_bus[1];
assign cfg_coladdrwidth[2] = hmc_inst_CFGCOLADDRWIDTH_bus[2];
assign cfg_coladdrwidth[3] = hmc_inst_CFGCOLADDRWIDTH_bus[3];
assign cfg_coladdrwidth[4] = hmc_inst_CFGCOLADDRWIDTH_bus[4];

assign cfg_csaddrwidth[0] = hmc_inst_CFGCSADDRWIDTH_bus[0];
assign cfg_csaddrwidth[1] = hmc_inst_CFGCSADDRWIDTH_bus[1];
assign cfg_csaddrwidth[2] = hmc_inst_CFGCSADDRWIDTH_bus[2];

assign cfg_devicewidth[0] = hmc_inst_CFGDEVICEWIDTH_bus[0];
assign cfg_devicewidth[1] = hmc_inst_CFGDEVICEWIDTH_bus[1];
assign cfg_devicewidth[2] = hmc_inst_CFGDEVICEWIDTH_bus[2];
assign cfg_devicewidth[3] = hmc_inst_CFGDEVICEWIDTH_bus[3];

assign cfg_interfacewidth[0] = hmc_inst_CFGINTERFACEWIDTH_bus[0];
assign cfg_interfacewidth[1] = hmc_inst_CFGINTERFACEWIDTH_bus[1];
assign cfg_interfacewidth[2] = hmc_inst_CFGINTERFACEWIDTH_bus[2];
assign cfg_interfacewidth[3] = hmc_inst_CFGINTERFACEWIDTH_bus[3];
assign cfg_interfacewidth[4] = hmc_inst_CFGINTERFACEWIDTH_bus[4];
assign cfg_interfacewidth[5] = hmc_inst_CFGINTERFACEWIDTH_bus[5];
assign cfg_interfacewidth[6] = hmc_inst_CFGINTERFACEWIDTH_bus[6];
assign cfg_interfacewidth[7] = hmc_inst_CFGINTERFACEWIDTH_bus[7];

assign cfg_rowaddrwidth[0] = hmc_inst_CFGROWADDRWIDTH_bus[0];
assign cfg_rowaddrwidth[1] = hmc_inst_CFGROWADDRWIDTH_bus[1];
assign cfg_rowaddrwidth[2] = hmc_inst_CFGROWADDRWIDTH_bus[2];
assign cfg_rowaddrwidth[3] = hmc_inst_CFGROWADDRWIDTH_bus[3];
assign cfg_rowaddrwidth[4] = hmc_inst_CFGROWADDRWIDTH_bus[4];

assign cfg_tcl[0] = hmc_inst_CFGTCL_bus[0];
assign cfg_tcl[1] = hmc_inst_CFGTCL_bus[1];
assign cfg_tcl[2] = hmc_inst_CFGTCL_bus[2];
assign cfg_tcl[3] = hmc_inst_CFGTCL_bus[3];
assign cfg_tcl[4] = hmc_inst_CFGTCL_bus[4];

assign cfg_tmrd[0] = hmc_inst_CFGTMRD_bus[0];
assign cfg_tmrd[1] = hmc_inst_CFGTMRD_bus[1];
assign cfg_tmrd[2] = hmc_inst_CFGTMRD_bus[2];
assign cfg_tmrd[3] = hmc_inst_CFGTMRD_bus[3];

assign cfg_trefi[0] = hmc_inst_CFGTREFI_bus[0];
assign cfg_trefi[1] = hmc_inst_CFGTREFI_bus[1];
assign cfg_trefi[2] = hmc_inst_CFGTREFI_bus[2];
assign cfg_trefi[3] = hmc_inst_CFGTREFI_bus[3];
assign cfg_trefi[4] = hmc_inst_CFGTREFI_bus[4];
assign cfg_trefi[5] = hmc_inst_CFGTREFI_bus[5];
assign cfg_trefi[6] = hmc_inst_CFGTREFI_bus[6];
assign cfg_trefi[7] = hmc_inst_CFGTREFI_bus[7];
assign cfg_trefi[8] = hmc_inst_CFGTREFI_bus[8];
assign cfg_trefi[9] = hmc_inst_CFGTREFI_bus[9];
assign cfg_trefi[10] = hmc_inst_CFGTREFI_bus[10];
assign cfg_trefi[11] = hmc_inst_CFGTREFI_bus[11];
assign cfg_trefi[12] = hmc_inst_CFGTREFI_bus[12];

assign cfg_trfc[0] = hmc_inst_CFGTRFC_bus[0];
assign cfg_trfc[1] = hmc_inst_CFGTRFC_bus[1];
assign cfg_trfc[2] = hmc_inst_CFGTRFC_bus[2];
assign cfg_trfc[3] = hmc_inst_CFGTRFC_bus[3];
assign cfg_trfc[4] = hmc_inst_CFGTRFC_bus[4];
assign cfg_trfc[5] = hmc_inst_CFGTRFC_bus[5];
assign cfg_trfc[6] = hmc_inst_CFGTRFC_bus[6];
assign cfg_trfc[7] = hmc_inst_CFGTRFC_bus[7];

assign cfg_twr[0] = hmc_inst_CFGTWR_bus[0];
assign cfg_twr[1] = hmc_inst_CFGTWR_bus[1];
assign cfg_twr[2] = hmc_inst_CFGTWR_bus[2];
assign cfg_twr[3] = hmc_inst_CFGTWR_bus[3];

assign afi_mem_clk_disable[0] = hmc_inst_CTLMEMCLKDISABLE_bus[0];

assign cfg_dramconfig[0] = hmc_inst_DRAMCONFIG_bus[0];
assign cfg_dramconfig[1] = hmc_inst_DRAMCONFIG_bus[1];
assign cfg_dramconfig[2] = hmc_inst_DRAMCONFIG_bus[2];
assign cfg_dramconfig[3] = hmc_inst_DRAMCONFIG_bus[3];
assign cfg_dramconfig[4] = hmc_inst_DRAMCONFIG_bus[4];
assign cfg_dramconfig[5] = hmc_inst_DRAMCONFIG_bus[5];
assign cfg_dramconfig[6] = hmc_inst_DRAMCONFIG_bus[6];
assign cfg_dramconfig[7] = hmc_inst_DRAMCONFIG_bus[7];
assign cfg_dramconfig[8] = hmc_inst_DRAMCONFIG_bus[8];
assign cfg_dramconfig[9] = hmc_inst_DRAMCONFIG_bus[9];
assign cfg_dramconfig[10] = hmc_inst_DRAMCONFIG_bus[10];
assign cfg_dramconfig[11] = hmc_inst_DRAMCONFIG_bus[11];
assign cfg_dramconfig[12] = hmc_inst_DRAMCONFIG_bus[12];
assign cfg_dramconfig[13] = hmc_inst_DRAMCONFIG_bus[13];
assign cfg_dramconfig[14] = hmc_inst_DRAMCONFIG_bus[14];
assign cfg_dramconfig[15] = hmc_inst_DRAMCONFIG_bus[15];
assign cfg_dramconfig[16] = hmc_inst_DRAMCONFIG_bus[16];
assign cfg_dramconfig[17] = hmc_inst_DRAMCONFIG_bus[17];
assign cfg_dramconfig[18] = hmc_inst_DRAMCONFIG_bus[18];
assign cfg_dramconfig[19] = hmc_inst_DRAMCONFIG_bus[19];
assign cfg_dramconfig[20] = hmc_inst_DRAMCONFIG_bus[20];

cyclonev_hmc hmc_inst(
	.afirdatavalid(afi_rdata_valid[0]),
	.csrclk(gnd),
	.csrdin(gnd),
	.csren(gnd),
	.ctlcalfail(afi_cal_fail),
	.ctlcalsuccess(afi_cal_success),
	.ctlclk(ctl_clk),
	.ctlresetn(ctl_reset_n),
	.globalresetn(gnd),
	.iavstcmdresetn0(vcc),
	.iavstcmdresetn1(vcc),
	.iavstcmdresetn2(vcc),
	.iavstcmdresetn3(vcc),
	.iavstcmdresetn4(vcc),
	.iavstcmdresetn5(vcc),
	.iavstrdclk0(gnd),
	.iavstrdclk1(gnd),
	.iavstrdclk2(gnd),
	.iavstrdclk3(gnd),
	.iavstrdready0(vcc),
	.iavstrdready1(vcc),
	.iavstrdready2(vcc),
	.iavstrdready3(vcc),
	.iavstrdresetn0(vcc),
	.iavstrdresetn1(vcc),
	.iavstrdresetn2(vcc),
	.iavstrdresetn3(vcc),
	.iavstwrackready0(vcc),
	.iavstwrackready1(vcc),
	.iavstwrackready2(vcc),
	.iavstwrackready3(vcc),
	.iavstwrackready4(vcc),
	.iavstwrackready5(vcc),
	.iavstwrclk0(gnd),
	.iavstwrclk1(gnd),
	.iavstwrclk2(gnd),
	.iavstwrclk3(gnd),
	.iavstwrresetn0(vcc),
	.iavstwrresetn1(vcc),
	.iavstwrresetn2(vcc),
	.iavstwrresetn3(vcc),
	.localdeeppowerdnreq(gnd),
	.localrefreshreq(gnd),
	.localselfrfshreq(gnd),
	.mmrbe(gnd),
	.mmrburstbegin(vcc),
	.mmrclk(gnd),
	.mmrreadreq(gnd),
	.mmrresetn(vcc),
	.mmrwritereq(gnd),
	.portclk0(gnd),
	.portclk1(gnd),
	.portclk2(gnd),
	.portclk3(gnd),
	.portclk4(gnd),
	.portclk5(gnd),
	.scanenable(gnd),
	.scbe(gnd),
	.scburstbegin(gnd),
	.scclk(gnd),
	.screadreq(gnd),
	.scresetn(vcc),
	.scwritereq(gnd),
	.afirdata({afi_rdata[79],afi_rdata[78],afi_rdata[77],afi_rdata[76],afi_rdata[75],afi_rdata[74],afi_rdata[73],afi_rdata[72],afi_rdata[71],afi_rdata[70],afi_rdata[69],afi_rdata[68],afi_rdata[67],afi_rdata[66],afi_rdata[65],afi_rdata[64],afi_rdata[63],afi_rdata[62],afi_rdata[61],afi_rdata[60],afi_rdata[59],afi_rdata[58],afi_rdata[57],afi_rdata[56],afi_rdata[55],afi_rdata[54],afi_rdata[53],afi_rdata[52],
afi_rdata[51],afi_rdata[50],afi_rdata[49],afi_rdata[48],afi_rdata[47],afi_rdata[46],afi_rdata[45],afi_rdata[44],afi_rdata[43],afi_rdata[42],afi_rdata[41],afi_rdata[40],afi_rdata[39],afi_rdata[38],afi_rdata[37],afi_rdata[36],afi_rdata[35],afi_rdata[34],afi_rdata[33],afi_rdata[32],afi_rdata[31],afi_rdata[30],afi_rdata[29],afi_rdata[28],afi_rdata[27],afi_rdata[26],afi_rdata[25],afi_rdata[24],
afi_rdata[23],afi_rdata[22],afi_rdata[21],afi_rdata[20],afi_rdata[19],afi_rdata[18],afi_rdata[17],afi_rdata[16],afi_rdata[15],afi_rdata[14],afi_rdata[13],afi_rdata[12],afi_rdata[11],afi_rdata[10],afi_rdata[9],afi_rdata[8],afi_rdata[7],afi_rdata[6],afi_rdata[5],afi_rdata[4],afi_rdata[3],afi_rdata[2],afi_rdata[1],afi_rdata[0]}),
	.afiseqbusy({gnd,gnd}),
	.afiwlat({afi_wlat[3],afi_wlat[2],afi_wlat[1],afi_wlat[0]}),
	.bondingin1({gnd,gnd,gnd,gnd}),
	.bondingin2({gnd,gnd,gnd,gnd,gnd,gnd}),
	.bondingin3({gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata4({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata5({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.localdeeppowerdnchip({gnd,gnd}),
	.localrefreshchip({gnd,gnd}),
	.localselfrfshchip({gnd,gnd}),
	.mmraddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.mmrburstcount({gnd,vcc}),
	.mmrwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scburstcount({gnd,gnd}),
	.scwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.aficasn(afi_cas_n[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.csrdout(),
	.ctlcalreq(),
	.ctlinitreq(),
	.localdeeppowerdnack(),
	.localinitdone(),
	.localpowerdownack(),
	.localrefreshack(),
	.localselfrfshack(),
	.localstsctlempty(),
	.mmrrdatavalid(),
	.mmrwaitrequest(),
	.oammready0(),
	.oammready1(),
	.oammready2(),
	.oammready3(),
	.oammready4(),
	.oammready5(),
	.ordavstvalid0(),
	.ordavstvalid1(),
	.ordavstvalid2(),
	.ordavstvalid3(),
	.owrackavstdata0(),
	.owrackavstdata1(),
	.owrackavstdata2(),
	.owrackavstdata3(),
	.owrackavstdata4(),
	.owrackavstdata5(),
	.owrackavstvalid0(),
	.owrackavstvalid1(),
	.owrackavstvalid2(),
	.owrackavstvalid3(),
	.owrackavstvalid4(),
	.owrackavstvalid5(),
	.scrdatavalid(),
	.scwaitrequest(),
	.afiaddr(hmc_inst_AFIADDR_bus),
	.afiba(hmc_inst_AFIBA_bus),
	.aficke(hmc_inst_AFICKE_bus),
	.aficsn(hmc_inst_AFICSN_bus),
	.afictllongidle(),
	.afictlrefreshdone(),
	.afidm(hmc_inst_AFIDM_bus),
	.afidqsburst(hmc_inst_AFIDQSBURST_bus),
	.afiodt(hmc_inst_AFIODT_bus),
	.afirdataen(hmc_inst_AFIRDATAEN_bus),
	.afirdataenfull(hmc_inst_AFIRDATAENFULL_bus),
	.afiwdata(hmc_inst_AFIWDATA_bus),
	.afiwdatavalid(hmc_inst_AFIWDATAVALID_bus),
	.bondingout1(),
	.bondingout2(),
	.bondingout3(),
	.cfgaddlat(hmc_inst_CFGADDLAT_bus),
	.cfgbankaddrwidth(hmc_inst_CFGBANKADDRWIDTH_bus),
	.cfgcaswrlat(hmc_inst_CFGCASWRLAT_bus),
	.cfgcoladdrwidth(hmc_inst_CFGCOLADDRWIDTH_bus),
	.cfgcsaddrwidth(hmc_inst_CFGCSADDRWIDTH_bus),
	.cfgdevicewidth(hmc_inst_CFGDEVICEWIDTH_bus),
	.cfginterfacewidth(hmc_inst_CFGINTERFACEWIDTH_bus),
	.cfgrowaddrwidth(hmc_inst_CFGROWADDRWIDTH_bus),
	.cfgtcl(hmc_inst_CFGTCL_bus),
	.cfgtmrd(hmc_inst_CFGTMRD_bus),
	.cfgtrefi(hmc_inst_CFGTREFI_bus),
	.cfgtrfc(hmc_inst_CFGTRFC_bus),
	.cfgtwr(hmc_inst_CFGTWR_bus),
	.ctlcalbytelaneseln(),
	.ctlmemclkdisable(hmc_inst_CTLMEMCLKDISABLE_bus),
	.dramconfig(hmc_inst_DRAMCONFIG_bus),
	.mmrrdata(),
	.ordavstdata0(),
	.ordavstdata1(),
	.ordavstdata2(),
	.ordavstdata3(),
	.scrdata());
defparam hmc_inst.attr_counter_one_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_reset = "disabled";
defparam hmc_inst.attr_counter_zero_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_reset = "disabled";
defparam hmc_inst.attr_debug_select_byte = 32'b00000000000000000000000000000000;
defparam hmc_inst.attr_static_config_valid = "disabled";
defparam hmc_inst.auto_pch_enable_0 = "disabled";
defparam hmc_inst.auto_pch_enable_1 = "disabled";
defparam hmc_inst.auto_pch_enable_2 = "disabled";
defparam hmc_inst.auto_pch_enable_3 = "disabled";
defparam hmc_inst.auto_pch_enable_4 = "disabled";
defparam hmc_inst.auto_pch_enable_5 = "disabled";
defparam hmc_inst.cal_req = "disabled";
defparam hmc_inst.cfg_burst_length = "bl_8";
defparam hmc_inst.cfg_interface_width = "dwidth_32";
defparam hmc_inst.cfg_self_rfsh_exit_cycles = "self_rfsh_exit_cycles_512";
defparam hmc_inst.cfg_starve_limit = "starve_limit_10";
defparam hmc_inst.cfg_type = "ddr3";
defparam hmc_inst.clr_intr = "no_clr_intr";
defparam hmc_inst.cmd_port_in_use_0 = "false";
defparam hmc_inst.cmd_port_in_use_1 = "false";
defparam hmc_inst.cmd_port_in_use_2 = "false";
defparam hmc_inst.cmd_port_in_use_3 = "false";
defparam hmc_inst.cmd_port_in_use_4 = "false";
defparam hmc_inst.cmd_port_in_use_5 = "false";
defparam hmc_inst.cport0_rdy_almost_full = "not_full";
defparam hmc_inst.cport0_rfifo_map = "fifo_0";
defparam hmc_inst.cport0_type = "disable";
defparam hmc_inst.cport0_wfifo_map = "fifo_0";
defparam hmc_inst.cport1_rdy_almost_full = "not_full";
defparam hmc_inst.cport1_rfifo_map = "fifo_0";
defparam hmc_inst.cport1_type = "disable";
defparam hmc_inst.cport1_wfifo_map = "fifo_0";
defparam hmc_inst.cport2_rdy_almost_full = "not_full";
defparam hmc_inst.cport2_rfifo_map = "fifo_0";
defparam hmc_inst.cport2_type = "disable";
defparam hmc_inst.cport2_wfifo_map = "fifo_0";
defparam hmc_inst.cport3_rdy_almost_full = "not_full";
defparam hmc_inst.cport3_rfifo_map = "fifo_0";
defparam hmc_inst.cport3_type = "disable";
defparam hmc_inst.cport3_wfifo_map = "fifo_0";
defparam hmc_inst.cport4_rdy_almost_full = "not_full";
defparam hmc_inst.cport4_rfifo_map = "fifo_0";
defparam hmc_inst.cport4_type = "disable";
defparam hmc_inst.cport4_wfifo_map = "fifo_0";
defparam hmc_inst.cport5_rdy_almost_full = "not_full";
defparam hmc_inst.cport5_rfifo_map = "fifo_0";
defparam hmc_inst.cport5_type = "disable";
defparam hmc_inst.cport5_wfifo_map = "fifo_0";
defparam hmc_inst.ctl_addr_order = "chip_row_bank_col";
defparam hmc_inst.ctl_ecc_enabled = "ctl_ecc_disabled";
defparam hmc_inst.ctl_ecc_rmw_enabled = "ctl_ecc_rmw_disabled";
defparam hmc_inst.ctl_regdimm_enabled = "regdimm_disabled";
defparam hmc_inst.ctl_usr_refresh = "ctl_usr_refresh_disabled";
defparam hmc_inst.ctrl_width = "data_width_64_bit";
defparam hmc_inst.cyc_to_rld_jars_0 = 1;
defparam hmc_inst.cyc_to_rld_jars_1 = 1;
defparam hmc_inst.cyc_to_rld_jars_2 = 1;
defparam hmc_inst.cyc_to_rld_jars_3 = 1;
defparam hmc_inst.cyc_to_rld_jars_4 = 1;
defparam hmc_inst.cyc_to_rld_jars_5 = 1;
defparam hmc_inst.delay_bonding = "bonding_latency_0";
defparam hmc_inst.dfx_bypass_enable = "dfx_bypass_disabled";
defparam hmc_inst.disable_merging = "merging_enabled";
defparam hmc_inst.ecc_dq_width = "ecc_dq_width_0";
defparam hmc_inst.enable_atpg = "disabled";
defparam hmc_inst.enable_bonding_0 = "disabled";
defparam hmc_inst.enable_bonding_1 = "disabled";
defparam hmc_inst.enable_bonding_2 = "disabled";
defparam hmc_inst.enable_bonding_3 = "disabled";
defparam hmc_inst.enable_bonding_4 = "disabled";
defparam hmc_inst.enable_bonding_5 = "disabled";
defparam hmc_inst.enable_bonding_wrapback = "disabled";
defparam hmc_inst.enable_burst_interrupt = "disabled";
defparam hmc_inst.enable_burst_terminate = "disabled";
defparam hmc_inst.enable_dqs_tracking = "enabled";
defparam hmc_inst.enable_ecc_code_overwrites = "disabled";
defparam hmc_inst.enable_fast_exit_ppd = "disabled";
defparam hmc_inst.enable_intr = "disabled";
defparam hmc_inst.enable_no_dm = "disabled";
defparam hmc_inst.enable_pipelineglobal = "disabled";
defparam hmc_inst.extra_ctl_clk_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_act_to_act_diff_bank = 0;
defparam hmc_inst.extra_ctl_clk_act_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_act_to_rdwr = 0;
defparam hmc_inst.extra_ctl_clk_arf_period = 0;
defparam hmc_inst.extra_ctl_clk_arf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_four_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_pch_all_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pch_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pdn_period = 0;
defparam hmc_inst.extra_ctl_clk_pdn_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd_diff_chip = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_wr = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_bc = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_diff_chip = 2;
defparam hmc_inst.extra_ctl_clk_srf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_srf_to_zq_cal = 0;
defparam hmc_inst.extra_ctl_clk_wr_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_rd = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_bc = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_diff_chip = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_wr = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_wr_diff_chip = 0;
defparam hmc_inst.gen_dbe = "gen_dbe_disabled";
defparam hmc_inst.gen_sbe = "gen_sbe_disabled";
defparam hmc_inst.inc_sync = "fifo_set_2";
defparam hmc_inst.local_if_cs_width = "addr_width_0";
defparam hmc_inst.mask_corr_dropped_intr = "disabled";
defparam hmc_inst.mask_dbe_intr = "disabled";
defparam hmc_inst.mask_sbe_intr = "disabled";
defparam hmc_inst.mem_auto_pd_cycles = 0;
defparam hmc_inst.mem_clk_entry_cycles = 10;
defparam hmc_inst.mem_if_al = "al_0";
defparam hmc_inst.mem_if_bankaddr_width = "addr_width_3";
defparam hmc_inst.mem_if_burstlength = "mem_if_burstlength_8";
defparam hmc_inst.mem_if_coladdr_width = "addr_width_10";
defparam hmc_inst.mem_if_cs_per_rank = "mem_if_cs_per_rank_1";
defparam hmc_inst.mem_if_cs_width = "mem_if_cs_width_1";
defparam hmc_inst.mem_if_dq_per_chip = "mem_if_dq_per_chip_8";
defparam hmc_inst.mem_if_dqs_width = "dqs_width_4";
defparam hmc_inst.mem_if_dwidth = "mem_if_dwidth_32";
defparam hmc_inst.mem_if_memtype = "ddr3_sdram";
defparam hmc_inst.mem_if_rowaddr_width = "addr_width_15";
defparam hmc_inst.mem_if_speedbin = "ddr3_1600_8_8_8";
defparam hmc_inst.mem_if_tccd = "tccd_4";
defparam hmc_inst.mem_if_tcl = "tcl_7";
defparam hmc_inst.mem_if_tcwl = "tcwl_7";
defparam hmc_inst.mem_if_tfaw = "tfaw_15";
defparam hmc_inst.mem_if_tmrd = "tmrd_4";
defparam hmc_inst.mem_if_tras = "tras_14";
defparam hmc_inst.mem_if_trc = "trc_20";
defparam hmc_inst.mem_if_trcd = "trcd_6";
defparam hmc_inst.mem_if_trefi = 3120;
defparam hmc_inst.mem_if_trfc = 120;
defparam hmc_inst.mem_if_trp = "trp_6";
defparam hmc_inst.mem_if_trrd = "trrd_3";
defparam hmc_inst.mem_if_trtp = "trtp_3";
defparam hmc_inst.mem_if_twr = "twr_6";
defparam hmc_inst.mem_if_twtr = "twtr_4";
defparam hmc_inst.mmr_cfg_mem_bl = "mp_bl_8";
defparam hmc_inst.output_regd = "disabled";
defparam hmc_inst.pdn_exit_cycles = "slow_exit";
defparam hmc_inst.port0_width = "port_32_bit";
defparam hmc_inst.port1_width = "port_32_bit";
defparam hmc_inst.port2_width = "port_32_bit";
defparam hmc_inst.port3_width = "port_32_bit";
defparam hmc_inst.port4_width = "port_32_bit";
defparam hmc_inst.port5_width = "port_32_bit";
defparam hmc_inst.power_saving_exit_cycles = 5;
defparam hmc_inst.priority_0_0 = "weight_0";
defparam hmc_inst.priority_0_1 = "weight_0";
defparam hmc_inst.priority_0_2 = "weight_0";
defparam hmc_inst.priority_0_3 = "weight_0";
defparam hmc_inst.priority_0_4 = "weight_0";
defparam hmc_inst.priority_0_5 = "weight_0";
defparam hmc_inst.priority_1_0 = "weight_0";
defparam hmc_inst.priority_1_1 = "weight_0";
defparam hmc_inst.priority_1_2 = "weight_0";
defparam hmc_inst.priority_1_3 = "weight_0";
defparam hmc_inst.priority_1_4 = "weight_0";
defparam hmc_inst.priority_1_5 = "weight_0";
defparam hmc_inst.priority_2_0 = "weight_0";
defparam hmc_inst.priority_2_1 = "weight_0";
defparam hmc_inst.priority_2_2 = "weight_0";
defparam hmc_inst.priority_2_3 = "weight_0";
defparam hmc_inst.priority_2_4 = "weight_0";
defparam hmc_inst.priority_2_5 = "weight_0";
defparam hmc_inst.priority_3_0 = "weight_0";
defparam hmc_inst.priority_3_1 = "weight_0";
defparam hmc_inst.priority_3_2 = "weight_0";
defparam hmc_inst.priority_3_3 = "weight_0";
defparam hmc_inst.priority_3_4 = "weight_0";
defparam hmc_inst.priority_3_5 = "weight_0";
defparam hmc_inst.priority_4_0 = "weight_0";
defparam hmc_inst.priority_4_1 = "weight_0";
defparam hmc_inst.priority_4_2 = "weight_0";
defparam hmc_inst.priority_4_3 = "weight_0";
defparam hmc_inst.priority_4_4 = "weight_0";
defparam hmc_inst.priority_4_5 = "weight_0";
defparam hmc_inst.priority_5_0 = "weight_0";
defparam hmc_inst.priority_5_1 = "weight_0";
defparam hmc_inst.priority_5_2 = "weight_0";
defparam hmc_inst.priority_5_3 = "weight_0";
defparam hmc_inst.priority_5_4 = "weight_0";
defparam hmc_inst.priority_5_5 = "weight_0";
defparam hmc_inst.priority_6_0 = "weight_0";
defparam hmc_inst.priority_6_1 = "weight_0";
defparam hmc_inst.priority_6_2 = "weight_0";
defparam hmc_inst.priority_6_3 = "weight_0";
defparam hmc_inst.priority_6_4 = "weight_0";
defparam hmc_inst.priority_6_5 = "weight_0";
defparam hmc_inst.priority_7_0 = "weight_0";
defparam hmc_inst.priority_7_1 = "weight_0";
defparam hmc_inst.priority_7_2 = "weight_0";
defparam hmc_inst.priority_7_3 = "weight_0";
defparam hmc_inst.priority_7_4 = "weight_0";
defparam hmc_inst.priority_7_5 = "weight_0";
defparam hmc_inst.priority_remap = 0;
defparam hmc_inst.rcfg_static_weight_0 = "weight_0";
defparam hmc_inst.rcfg_static_weight_1 = "weight_0";
defparam hmc_inst.rcfg_static_weight_2 = "weight_0";
defparam hmc_inst.rcfg_static_weight_3 = "weight_0";
defparam hmc_inst.rcfg_static_weight_4 = "weight_0";
defparam hmc_inst.rcfg_static_weight_5 = "weight_0";
defparam hmc_inst.rcfg_sum_wt_priority_0 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_1 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_2 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_3 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_4 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_5 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_6 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_7 = 0;
defparam hmc_inst.rcfg_user_priority_0 = "priority_1";
defparam hmc_inst.rcfg_user_priority_1 = "priority_1";
defparam hmc_inst.rcfg_user_priority_2 = "priority_1";
defparam hmc_inst.rcfg_user_priority_3 = "priority_1";
defparam hmc_inst.rcfg_user_priority_4 = "priority_1";
defparam hmc_inst.rcfg_user_priority_5 = "priority_1";
defparam hmc_inst.rd_dwidth_0 = "dwidth_0";
defparam hmc_inst.rd_dwidth_1 = "dwidth_0";
defparam hmc_inst.rd_dwidth_2 = "dwidth_0";
defparam hmc_inst.rd_dwidth_3 = "dwidth_0";
defparam hmc_inst.rd_dwidth_4 = "dwidth_0";
defparam hmc_inst.rd_dwidth_5 = "dwidth_0";
defparam hmc_inst.rd_fifo_in_use_0 = "false";
defparam hmc_inst.rd_fifo_in_use_1 = "false";
defparam hmc_inst.rd_fifo_in_use_2 = "false";
defparam hmc_inst.rd_fifo_in_use_3 = "false";
defparam hmc_inst.rd_port_info_0 = "use_no";
defparam hmc_inst.rd_port_info_1 = "use_no";
defparam hmc_inst.rd_port_info_2 = "use_no";
defparam hmc_inst.rd_port_info_3 = "use_no";
defparam hmc_inst.rd_port_info_4 = "use_no";
defparam hmc_inst.rd_port_info_5 = "use_no";
defparam hmc_inst.read_odt_chip = "odt_disabled";
defparam hmc_inst.reorder_data = "data_reordering";
defparam hmc_inst.rfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.single_ready_0 = "concatenate_rdy";
defparam hmc_inst.single_ready_1 = "concatenate_rdy";
defparam hmc_inst.single_ready_2 = "concatenate_rdy";
defparam hmc_inst.single_ready_3 = "concatenate_rdy";
defparam hmc_inst.static_weight_0 = "weight_0";
defparam hmc_inst.static_weight_1 = "weight_0";
defparam hmc_inst.static_weight_2 = "weight_0";
defparam hmc_inst.static_weight_3 = "weight_0";
defparam hmc_inst.static_weight_4 = "weight_0";
defparam hmc_inst.static_weight_5 = "weight_0";
defparam hmc_inst.sum_wt_priority_0 = 0;
defparam hmc_inst.sum_wt_priority_1 = 0;
defparam hmc_inst.sum_wt_priority_2 = 0;
defparam hmc_inst.sum_wt_priority_3 = 0;
defparam hmc_inst.sum_wt_priority_4 = 0;
defparam hmc_inst.sum_wt_priority_5 = 0;
defparam hmc_inst.sum_wt_priority_6 = 0;
defparam hmc_inst.sum_wt_priority_7 = 0;
defparam hmc_inst.sync_mode_0 = "asynchronous";
defparam hmc_inst.sync_mode_1 = "asynchronous";
defparam hmc_inst.sync_mode_2 = "asynchronous";
defparam hmc_inst.sync_mode_3 = "asynchronous";
defparam hmc_inst.sync_mode_4 = "asynchronous";
defparam hmc_inst.sync_mode_5 = "asynchronous";
defparam hmc_inst.test_mode = "normal_mode";
defparam hmc_inst.thld_jar1_0 = "threshold_32";
defparam hmc_inst.thld_jar1_1 = "threshold_32";
defparam hmc_inst.thld_jar1_2 = "threshold_32";
defparam hmc_inst.thld_jar1_3 = "threshold_32";
defparam hmc_inst.thld_jar1_4 = "threshold_32";
defparam hmc_inst.thld_jar1_5 = "threshold_32";
defparam hmc_inst.thld_jar2_0 = "threshold_16";
defparam hmc_inst.thld_jar2_1 = "threshold_16";
defparam hmc_inst.thld_jar2_2 = "threshold_16";
defparam hmc_inst.thld_jar2_3 = "threshold_16";
defparam hmc_inst.thld_jar2_4 = "threshold_16";
defparam hmc_inst.thld_jar2_5 = "threshold_16";
defparam hmc_inst.use_almost_empty_0 = "empty";
defparam hmc_inst.use_almost_empty_1 = "empty";
defparam hmc_inst.use_almost_empty_2 = "empty";
defparam hmc_inst.use_almost_empty_3 = "empty";
defparam hmc_inst.user_ecc_en = "disable";
defparam hmc_inst.user_priority_0 = "priority_1";
defparam hmc_inst.user_priority_1 = "priority_1";
defparam hmc_inst.user_priority_2 = "priority_1";
defparam hmc_inst.user_priority_3 = "priority_1";
defparam hmc_inst.user_priority_4 = "priority_1";
defparam hmc_inst.user_priority_5 = "priority_1";
defparam hmc_inst.wfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo0_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo1_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo2_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo3_rdy_almost_full = "not_full";
defparam hmc_inst.wr_dwidth_0 = "dwidth_0";
defparam hmc_inst.wr_dwidth_1 = "dwidth_0";
defparam hmc_inst.wr_dwidth_2 = "dwidth_0";
defparam hmc_inst.wr_dwidth_3 = "dwidth_0";
defparam hmc_inst.wr_dwidth_4 = "dwidth_0";
defparam hmc_inst.wr_dwidth_5 = "dwidth_0";
defparam hmc_inst.wr_fifo_in_use_0 = "false";
defparam hmc_inst.wr_fifo_in_use_1 = "false";
defparam hmc_inst.wr_fifo_in_use_2 = "false";
defparam hmc_inst.wr_fifo_in_use_3 = "false";
defparam hmc_inst.wr_port_info_0 = "use_no";
defparam hmc_inst.wr_port_info_1 = "use_no";
defparam hmc_inst.wr_port_info_2 = "use_no";
defparam hmc_inst.wr_port_info_3 = "use_no";
defparam hmc_inst.wr_port_info_4 = "use_no";
defparam hmc_inst.wr_port_info_5 = "use_no";
defparam hmc_inst.write_odt_chip = "write_chip0_odt0_chip1";

endmodule

module soc_system_altera_mem_if_oct_cyclonev (
	parallelterminationcontrol,
	seriesterminationcontrol,
	oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[15:0] parallelterminationcontrol;
output 	[15:0] seriesterminationcontrol;
input 	oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sd1a_0~O_CLKUSRDFTOUT ;
wire \wire_sd1a_serdataout[0] ;

wire [15:0] sd2a_0_PARALLELTERMINATIONCONTROL_bus;
wire [15:0] sd2a_0_SERIESTERMINATIONCONTROL_bus;

assign parallelterminationcontrol[0] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[0];
assign parallelterminationcontrol[1] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[1];
assign parallelterminationcontrol[2] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[2];
assign parallelterminationcontrol[3] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[3];
assign parallelterminationcontrol[4] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[4];
assign parallelterminationcontrol[5] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[5];
assign parallelterminationcontrol[6] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[6];
assign parallelterminationcontrol[7] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[7];
assign parallelterminationcontrol[8] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[8];
assign parallelterminationcontrol[9] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[9];
assign parallelterminationcontrol[10] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[10];
assign parallelterminationcontrol[11] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[11];
assign parallelterminationcontrol[12] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[12];
assign parallelterminationcontrol[13] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[13];
assign parallelterminationcontrol[14] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[14];
assign parallelterminationcontrol[15] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[15];

assign seriesterminationcontrol[0] = sd2a_0_SERIESTERMINATIONCONTROL_bus[0];
assign seriesterminationcontrol[1] = sd2a_0_SERIESTERMINATIONCONTROL_bus[1];
assign seriesterminationcontrol[2] = sd2a_0_SERIESTERMINATIONCONTROL_bus[2];
assign seriesterminationcontrol[3] = sd2a_0_SERIESTERMINATIONCONTROL_bus[3];
assign seriesterminationcontrol[4] = sd2a_0_SERIESTERMINATIONCONTROL_bus[4];
assign seriesterminationcontrol[5] = sd2a_0_SERIESTERMINATIONCONTROL_bus[5];
assign seriesterminationcontrol[6] = sd2a_0_SERIESTERMINATIONCONTROL_bus[6];
assign seriesterminationcontrol[7] = sd2a_0_SERIESTERMINATIONCONTROL_bus[7];
assign seriesterminationcontrol[8] = sd2a_0_SERIESTERMINATIONCONTROL_bus[8];
assign seriesterminationcontrol[9] = sd2a_0_SERIESTERMINATIONCONTROL_bus[9];
assign seriesterminationcontrol[10] = sd2a_0_SERIESTERMINATIONCONTROL_bus[10];
assign seriesterminationcontrol[11] = sd2a_0_SERIESTERMINATIONCONTROL_bus[11];
assign seriesterminationcontrol[12] = sd2a_0_SERIESTERMINATIONCONTROL_bus[12];
assign seriesterminationcontrol[13] = sd2a_0_SERIESTERMINATIONCONTROL_bus[13];
assign seriesterminationcontrol[14] = sd2a_0_SERIESTERMINATIONCONTROL_bus[14];
assign seriesterminationcontrol[15] = sd2a_0_SERIESTERMINATIONCONTROL_bus[15];

cyclonev_termination_logic sd2a_0(
	.s2pload(gnd),
	.scanclk(gnd),
	.scanenable(gnd),
	.serdata(\wire_sd1a_serdataout[0] ),
	.enser(4'b0000),
	.parallelterminationcontrol(sd2a_0_PARALLELTERMINATIONCONTROL_bus),
	.seriesterminationcontrol(sd2a_0_SERIESTERMINATIONCONTROL_bus));

cyclonev_termination sd1a_0(
	.clkenusr(gnd),
	.clkusr(gnd),
	.enserusr(gnd),
	.nclrusr(gnd),
	.rzqin(oct_rzqin),
	.scanclk(gnd),
	.scanen(gnd),
	.scanin(gnd),
	.serdatafromcore(gnd),
	.serdatain(gnd),
	.otherenser(10'b0000000000),
	.clkusrdftout(\sd1a_0~O_CLKUSRDFTOUT ),
	.compoutrdn(),
	.compoutrup(),
	.enserout(),
	.scanout(),
	.serdataout(\wire_sd1a_serdataout[0] ),
	.serdatatocore());

endmodule

module soc_system_hps_sdram_p0 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid_0,
	ctl_reset_n,
	afi_rdata_0,
	afi_rdata_1,
	afi_rdata_2,
	afi_rdata_3,
	afi_rdata_4,
	afi_rdata_5,
	afi_rdata_6,
	afi_rdata_7,
	afi_rdata_8,
	afi_rdata_9,
	afi_rdata_10,
	afi_rdata_11,
	afi_rdata_12,
	afi_rdata_13,
	afi_rdata_14,
	afi_rdata_15,
	afi_rdata_16,
	afi_rdata_17,
	afi_rdata_18,
	afi_rdata_19,
	afi_rdata_20,
	afi_rdata_21,
	afi_rdata_22,
	afi_rdata_23,
	afi_rdata_24,
	afi_rdata_25,
	afi_rdata_26,
	afi_rdata_27,
	afi_rdata_28,
	afi_rdata_29,
	afi_rdata_30,
	afi_rdata_31,
	afi_rdata_32,
	afi_rdata_33,
	afi_rdata_34,
	afi_rdata_35,
	afi_rdata_36,
	afi_rdata_37,
	afi_rdata_38,
	afi_rdata_39,
	afi_rdata_40,
	afi_rdata_41,
	afi_rdata_42,
	afi_rdata_43,
	afi_rdata_44,
	afi_rdata_45,
	afi_rdata_46,
	afi_rdata_47,
	afi_rdata_48,
	afi_rdata_49,
	afi_rdata_50,
	afi_rdata_51,
	afi_rdata_52,
	afi_rdata_53,
	afi_rdata_54,
	afi_rdata_55,
	afi_rdata_56,
	afi_rdata_57,
	afi_rdata_58,
	afi_rdata_59,
	afi_rdata_60,
	afi_rdata_61,
	afi_rdata_62,
	afi_rdata_63,
	afi_rdata_64,
	afi_rdata_65,
	afi_rdata_66,
	afi_rdata_67,
	afi_rdata_68,
	afi_rdata_69,
	afi_rdata_70,
	afi_rdata_71,
	afi_rdata_72,
	afi_rdata_73,
	afi_rdata_74,
	afi_rdata_75,
	afi_rdata_76,
	afi_rdata_77,
	afi_rdata_78,
	afi_rdata_79,
	afi_wlat_0,
	afi_wlat_1,
	afi_wlat_2,
	afi_wlat_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n_0,
	afi_ras_n_0,
	afi_rst_n_0,
	afi_we_n_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_addr_14,
	afi_addr_15,
	afi_addr_16,
	afi_addr_17,
	afi_addr_18,
	afi_addr_19,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_cke_0,
	afi_cke_1,
	afi_cs_n_0,
	afi_cs_n_1,
	afi_dm_int_0,
	afi_dm_int_1,
	afi_dm_int_2,
	afi_dm_int_3,
	afi_dm_int_4,
	afi_dm_int_5,
	afi_dm_int_6,
	afi_dm_int_7,
	afi_dm_int_8,
	afi_dm_int_9,
	afi_dqs_burst_0,
	afi_dqs_burst_1,
	afi_dqs_burst_2,
	afi_dqs_burst_3,
	afi_dqs_burst_4,
	afi_odt_0,
	afi_odt_1,
	afi_rdata_en_0,
	afi_rdata_en_1,
	afi_rdata_en_2,
	afi_rdata_en_3,
	afi_rdata_en_4,
	afi_rdata_en_full_0,
	afi_rdata_en_full_1,
	afi_rdata_en_full_2,
	afi_rdata_en_full_3,
	afi_rdata_en_full_4,
	afi_wdata_int_0,
	afi_wdata_int_1,
	afi_wdata_int_2,
	afi_wdata_int_3,
	afi_wdata_int_4,
	afi_wdata_int_5,
	afi_wdata_int_6,
	afi_wdata_int_7,
	afi_wdata_int_8,
	afi_wdata_int_9,
	afi_wdata_int_10,
	afi_wdata_int_11,
	afi_wdata_int_12,
	afi_wdata_int_13,
	afi_wdata_int_14,
	afi_wdata_int_15,
	afi_wdata_int_16,
	afi_wdata_int_17,
	afi_wdata_int_18,
	afi_wdata_int_19,
	afi_wdata_int_20,
	afi_wdata_int_21,
	afi_wdata_int_22,
	afi_wdata_int_23,
	afi_wdata_int_24,
	afi_wdata_int_25,
	afi_wdata_int_26,
	afi_wdata_int_27,
	afi_wdata_int_28,
	afi_wdata_int_29,
	afi_wdata_int_30,
	afi_wdata_int_31,
	afi_wdata_int_32,
	afi_wdata_int_33,
	afi_wdata_int_34,
	afi_wdata_int_35,
	afi_wdata_int_36,
	afi_wdata_int_37,
	afi_wdata_int_38,
	afi_wdata_int_39,
	afi_wdata_int_40,
	afi_wdata_int_41,
	afi_wdata_int_42,
	afi_wdata_int_43,
	afi_wdata_int_44,
	afi_wdata_int_45,
	afi_wdata_int_46,
	afi_wdata_int_47,
	afi_wdata_int_48,
	afi_wdata_int_49,
	afi_wdata_int_50,
	afi_wdata_int_51,
	afi_wdata_int_52,
	afi_wdata_int_53,
	afi_wdata_int_54,
	afi_wdata_int_55,
	afi_wdata_int_56,
	afi_wdata_int_57,
	afi_wdata_int_58,
	afi_wdata_int_59,
	afi_wdata_int_60,
	afi_wdata_int_61,
	afi_wdata_int_62,
	afi_wdata_int_63,
	afi_wdata_int_64,
	afi_wdata_int_65,
	afi_wdata_int_66,
	afi_wdata_int_67,
	afi_wdata_int_68,
	afi_wdata_int_69,
	afi_wdata_int_70,
	afi_wdata_int_71,
	afi_wdata_int_72,
	afi_wdata_int_73,
	afi_wdata_int_74,
	afi_wdata_int_75,
	afi_wdata_int_76,
	afi_wdata_int_77,
	afi_wdata_int_78,
	afi_wdata_int_79,
	afi_wdata_valid_0,
	afi_wdata_valid_1,
	afi_wdata_valid_2,
	afi_wdata_valid_3,
	afi_wdata_valid_4,
	cfg_addlat_wire_0,
	cfg_addlat_wire_1,
	cfg_addlat_wire_2,
	cfg_addlat_wire_3,
	cfg_addlat_wire_4,
	cfg_bankaddrwidth_wire_0,
	cfg_bankaddrwidth_wire_1,
	cfg_bankaddrwidth_wire_2,
	cfg_caswrlat_wire_0,
	cfg_caswrlat_wire_1,
	cfg_caswrlat_wire_2,
	cfg_caswrlat_wire_3,
	cfg_coladdrwidth_wire_0,
	cfg_coladdrwidth_wire_1,
	cfg_coladdrwidth_wire_2,
	cfg_coladdrwidth_wire_3,
	cfg_coladdrwidth_wire_4,
	cfg_csaddrwidth_wire_0,
	cfg_csaddrwidth_wire_1,
	cfg_csaddrwidth_wire_2,
	cfg_devicewidth_wire_0,
	cfg_devicewidth_wire_1,
	cfg_devicewidth_wire_2,
	cfg_devicewidth_wire_3,
	cfg_interfacewidth_wire_0,
	cfg_interfacewidth_wire_1,
	cfg_interfacewidth_wire_2,
	cfg_interfacewidth_wire_3,
	cfg_interfacewidth_wire_4,
	cfg_interfacewidth_wire_5,
	cfg_interfacewidth_wire_6,
	cfg_interfacewidth_wire_7,
	cfg_rowaddrwidth_wire_0,
	cfg_rowaddrwidth_wire_1,
	cfg_rowaddrwidth_wire_2,
	cfg_rowaddrwidth_wire_3,
	cfg_rowaddrwidth_wire_4,
	cfg_tcl_wire_0,
	cfg_tcl_wire_1,
	cfg_tcl_wire_2,
	cfg_tcl_wire_3,
	cfg_tcl_wire_4,
	cfg_tmrd_wire_0,
	cfg_tmrd_wire_1,
	cfg_tmrd_wire_2,
	cfg_tmrd_wire_3,
	cfg_trefi_wire_0,
	cfg_trefi_wire_1,
	cfg_trefi_wire_2,
	cfg_trefi_wire_3,
	cfg_trefi_wire_4,
	cfg_trefi_wire_5,
	cfg_trefi_wire_6,
	cfg_trefi_wire_7,
	cfg_trefi_wire_8,
	cfg_trefi_wire_9,
	cfg_trefi_wire_10,
	cfg_trefi_wire_11,
	cfg_trefi_wire_12,
	cfg_trfc_wire_0,
	cfg_trfc_wire_1,
	cfg_trfc_wire_2,
	cfg_trfc_wire_3,
	cfg_trfc_wire_4,
	cfg_trfc_wire_5,
	cfg_trfc_wire_6,
	cfg_trfc_wire_7,
	cfg_twr_wire_0,
	cfg_twr_wire_1,
	cfg_twr_wire_2,
	cfg_twr_wire_3,
	afi_mem_clk_disable_0,
	cfg_dramconfig_wire_0,
	cfg_dramconfig_wire_1,
	cfg_dramconfig_wire_2,
	cfg_dramconfig_wire_3,
	cfg_dramconfig_wire_4,
	cfg_dramconfig_wire_5,
	cfg_dramconfig_wire_6,
	cfg_dramconfig_wire_7,
	cfg_dramconfig_wire_8,
	cfg_dramconfig_wire_9,
	cfg_dramconfig_wire_10,
	cfg_dramconfig_wire_11,
	cfg_dramconfig_wire_12,
	cfg_dramconfig_wire_13,
	cfg_dramconfig_wire_14,
	cfg_dramconfig_wire_15,
	cfg_dramconfig_wire_16,
	cfg_dramconfig_wire_17,
	cfg_dramconfig_wire_18,
	cfg_dramconfig_wire_19,
	cfg_dramconfig_wire_20,
	leveled_dqs_clocks_0,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	afi_rdata_valid_0;
output 	ctl_reset_n;
output 	afi_rdata_0;
output 	afi_rdata_1;
output 	afi_rdata_2;
output 	afi_rdata_3;
output 	afi_rdata_4;
output 	afi_rdata_5;
output 	afi_rdata_6;
output 	afi_rdata_7;
output 	afi_rdata_8;
output 	afi_rdata_9;
output 	afi_rdata_10;
output 	afi_rdata_11;
output 	afi_rdata_12;
output 	afi_rdata_13;
output 	afi_rdata_14;
output 	afi_rdata_15;
output 	afi_rdata_16;
output 	afi_rdata_17;
output 	afi_rdata_18;
output 	afi_rdata_19;
output 	afi_rdata_20;
output 	afi_rdata_21;
output 	afi_rdata_22;
output 	afi_rdata_23;
output 	afi_rdata_24;
output 	afi_rdata_25;
output 	afi_rdata_26;
output 	afi_rdata_27;
output 	afi_rdata_28;
output 	afi_rdata_29;
output 	afi_rdata_30;
output 	afi_rdata_31;
output 	afi_rdata_32;
output 	afi_rdata_33;
output 	afi_rdata_34;
output 	afi_rdata_35;
output 	afi_rdata_36;
output 	afi_rdata_37;
output 	afi_rdata_38;
output 	afi_rdata_39;
output 	afi_rdata_40;
output 	afi_rdata_41;
output 	afi_rdata_42;
output 	afi_rdata_43;
output 	afi_rdata_44;
output 	afi_rdata_45;
output 	afi_rdata_46;
output 	afi_rdata_47;
output 	afi_rdata_48;
output 	afi_rdata_49;
output 	afi_rdata_50;
output 	afi_rdata_51;
output 	afi_rdata_52;
output 	afi_rdata_53;
output 	afi_rdata_54;
output 	afi_rdata_55;
output 	afi_rdata_56;
output 	afi_rdata_57;
output 	afi_rdata_58;
output 	afi_rdata_59;
output 	afi_rdata_60;
output 	afi_rdata_61;
output 	afi_rdata_62;
output 	afi_rdata_63;
output 	afi_rdata_64;
output 	afi_rdata_65;
output 	afi_rdata_66;
output 	afi_rdata_67;
output 	afi_rdata_68;
output 	afi_rdata_69;
output 	afi_rdata_70;
output 	afi_rdata_71;
output 	afi_rdata_72;
output 	afi_rdata_73;
output 	afi_rdata_74;
output 	afi_rdata_75;
output 	afi_rdata_76;
output 	afi_rdata_77;
output 	afi_rdata_78;
output 	afi_rdata_79;
output 	afi_wlat_0;
output 	afi_wlat_1;
output 	afi_wlat_2;
output 	afi_wlat_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	afi_cas_n_0;
input 	afi_ras_n_0;
input 	afi_rst_n_0;
input 	afi_we_n_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_addr_14;
input 	afi_addr_15;
input 	afi_addr_16;
input 	afi_addr_17;
input 	afi_addr_18;
input 	afi_addr_19;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_cke_0;
input 	afi_cke_1;
input 	afi_cs_n_0;
input 	afi_cs_n_1;
input 	afi_dm_int_0;
input 	afi_dm_int_1;
input 	afi_dm_int_2;
input 	afi_dm_int_3;
input 	afi_dm_int_4;
input 	afi_dm_int_5;
input 	afi_dm_int_6;
input 	afi_dm_int_7;
input 	afi_dm_int_8;
input 	afi_dm_int_9;
input 	afi_dqs_burst_0;
input 	afi_dqs_burst_1;
input 	afi_dqs_burst_2;
input 	afi_dqs_burst_3;
input 	afi_dqs_burst_4;
input 	afi_odt_0;
input 	afi_odt_1;
input 	afi_rdata_en_0;
input 	afi_rdata_en_1;
input 	afi_rdata_en_2;
input 	afi_rdata_en_3;
input 	afi_rdata_en_4;
input 	afi_rdata_en_full_0;
input 	afi_rdata_en_full_1;
input 	afi_rdata_en_full_2;
input 	afi_rdata_en_full_3;
input 	afi_rdata_en_full_4;
input 	afi_wdata_int_0;
input 	afi_wdata_int_1;
input 	afi_wdata_int_2;
input 	afi_wdata_int_3;
input 	afi_wdata_int_4;
input 	afi_wdata_int_5;
input 	afi_wdata_int_6;
input 	afi_wdata_int_7;
input 	afi_wdata_int_8;
input 	afi_wdata_int_9;
input 	afi_wdata_int_10;
input 	afi_wdata_int_11;
input 	afi_wdata_int_12;
input 	afi_wdata_int_13;
input 	afi_wdata_int_14;
input 	afi_wdata_int_15;
input 	afi_wdata_int_16;
input 	afi_wdata_int_17;
input 	afi_wdata_int_18;
input 	afi_wdata_int_19;
input 	afi_wdata_int_20;
input 	afi_wdata_int_21;
input 	afi_wdata_int_22;
input 	afi_wdata_int_23;
input 	afi_wdata_int_24;
input 	afi_wdata_int_25;
input 	afi_wdata_int_26;
input 	afi_wdata_int_27;
input 	afi_wdata_int_28;
input 	afi_wdata_int_29;
input 	afi_wdata_int_30;
input 	afi_wdata_int_31;
input 	afi_wdata_int_32;
input 	afi_wdata_int_33;
input 	afi_wdata_int_34;
input 	afi_wdata_int_35;
input 	afi_wdata_int_36;
input 	afi_wdata_int_37;
input 	afi_wdata_int_38;
input 	afi_wdata_int_39;
input 	afi_wdata_int_40;
input 	afi_wdata_int_41;
input 	afi_wdata_int_42;
input 	afi_wdata_int_43;
input 	afi_wdata_int_44;
input 	afi_wdata_int_45;
input 	afi_wdata_int_46;
input 	afi_wdata_int_47;
input 	afi_wdata_int_48;
input 	afi_wdata_int_49;
input 	afi_wdata_int_50;
input 	afi_wdata_int_51;
input 	afi_wdata_int_52;
input 	afi_wdata_int_53;
input 	afi_wdata_int_54;
input 	afi_wdata_int_55;
input 	afi_wdata_int_56;
input 	afi_wdata_int_57;
input 	afi_wdata_int_58;
input 	afi_wdata_int_59;
input 	afi_wdata_int_60;
input 	afi_wdata_int_61;
input 	afi_wdata_int_62;
input 	afi_wdata_int_63;
input 	afi_wdata_int_64;
input 	afi_wdata_int_65;
input 	afi_wdata_int_66;
input 	afi_wdata_int_67;
input 	afi_wdata_int_68;
input 	afi_wdata_int_69;
input 	afi_wdata_int_70;
input 	afi_wdata_int_71;
input 	afi_wdata_int_72;
input 	afi_wdata_int_73;
input 	afi_wdata_int_74;
input 	afi_wdata_int_75;
input 	afi_wdata_int_76;
input 	afi_wdata_int_77;
input 	afi_wdata_int_78;
input 	afi_wdata_int_79;
input 	afi_wdata_valid_0;
input 	afi_wdata_valid_1;
input 	afi_wdata_valid_2;
input 	afi_wdata_valid_3;
input 	afi_wdata_valid_4;
input 	cfg_addlat_wire_0;
input 	cfg_addlat_wire_1;
input 	cfg_addlat_wire_2;
input 	cfg_addlat_wire_3;
input 	cfg_addlat_wire_4;
input 	cfg_bankaddrwidth_wire_0;
input 	cfg_bankaddrwidth_wire_1;
input 	cfg_bankaddrwidth_wire_2;
input 	cfg_caswrlat_wire_0;
input 	cfg_caswrlat_wire_1;
input 	cfg_caswrlat_wire_2;
input 	cfg_caswrlat_wire_3;
input 	cfg_coladdrwidth_wire_0;
input 	cfg_coladdrwidth_wire_1;
input 	cfg_coladdrwidth_wire_2;
input 	cfg_coladdrwidth_wire_3;
input 	cfg_coladdrwidth_wire_4;
input 	cfg_csaddrwidth_wire_0;
input 	cfg_csaddrwidth_wire_1;
input 	cfg_csaddrwidth_wire_2;
input 	cfg_devicewidth_wire_0;
input 	cfg_devicewidth_wire_1;
input 	cfg_devicewidth_wire_2;
input 	cfg_devicewidth_wire_3;
input 	cfg_interfacewidth_wire_0;
input 	cfg_interfacewidth_wire_1;
input 	cfg_interfacewidth_wire_2;
input 	cfg_interfacewidth_wire_3;
input 	cfg_interfacewidth_wire_4;
input 	cfg_interfacewidth_wire_5;
input 	cfg_interfacewidth_wire_6;
input 	cfg_interfacewidth_wire_7;
input 	cfg_rowaddrwidth_wire_0;
input 	cfg_rowaddrwidth_wire_1;
input 	cfg_rowaddrwidth_wire_2;
input 	cfg_rowaddrwidth_wire_3;
input 	cfg_rowaddrwidth_wire_4;
input 	cfg_tcl_wire_0;
input 	cfg_tcl_wire_1;
input 	cfg_tcl_wire_2;
input 	cfg_tcl_wire_3;
input 	cfg_tcl_wire_4;
input 	cfg_tmrd_wire_0;
input 	cfg_tmrd_wire_1;
input 	cfg_tmrd_wire_2;
input 	cfg_tmrd_wire_3;
input 	cfg_trefi_wire_0;
input 	cfg_trefi_wire_1;
input 	cfg_trefi_wire_2;
input 	cfg_trefi_wire_3;
input 	cfg_trefi_wire_4;
input 	cfg_trefi_wire_5;
input 	cfg_trefi_wire_6;
input 	cfg_trefi_wire_7;
input 	cfg_trefi_wire_8;
input 	cfg_trefi_wire_9;
input 	cfg_trefi_wire_10;
input 	cfg_trefi_wire_11;
input 	cfg_trefi_wire_12;
input 	cfg_trfc_wire_0;
input 	cfg_trfc_wire_1;
input 	cfg_trfc_wire_2;
input 	cfg_trfc_wire_3;
input 	cfg_trfc_wire_4;
input 	cfg_trfc_wire_5;
input 	cfg_trfc_wire_6;
input 	cfg_trfc_wire_7;
input 	cfg_twr_wire_0;
input 	cfg_twr_wire_1;
input 	cfg_twr_wire_2;
input 	cfg_twr_wire_3;
input 	afi_mem_clk_disable_0;
input 	cfg_dramconfig_wire_0;
input 	cfg_dramconfig_wire_1;
input 	cfg_dramconfig_wire_2;
input 	cfg_dramconfig_wire_3;
input 	cfg_dramconfig_wire_4;
input 	cfg_dramconfig_wire_5;
input 	cfg_dramconfig_wire_6;
input 	cfg_dramconfig_wire_7;
input 	cfg_dramconfig_wire_8;
input 	cfg_dramconfig_wire_9;
input 	cfg_dramconfig_wire_10;
input 	cfg_dramconfig_wire_11;
input 	cfg_dramconfig_wire_12;
input 	cfg_dramconfig_wire_13;
input 	cfg_dramconfig_wire_14;
input 	cfg_dramconfig_wire_15;
input 	cfg_dramconfig_wire_16;
input 	cfg_dramconfig_wire_17;
input 	cfg_dramconfig_wire_18;
input 	cfg_dramconfig_wire_19;
input 	cfg_dramconfig_wire_20;
output 	leveled_dqs_clocks_0;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_hps_sdram_p0_acv_hard_memphy umemphy(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(afi_cal_fail),
	.afi_cal_success(afi_cal_success),
	.afi_rdata_valid({afi_rdata_valid_0}),
	.ctl_reset_n(ctl_reset_n),
	.afi_rdata({afi_rdata_79,afi_rdata_78,afi_rdata_77,afi_rdata_76,afi_rdata_75,afi_rdata_74,afi_rdata_73,afi_rdata_72,afi_rdata_71,afi_rdata_70,afi_rdata_69,afi_rdata_68,afi_rdata_67,afi_rdata_66,afi_rdata_65,afi_rdata_64,afi_rdata_63,afi_rdata_62,afi_rdata_61,afi_rdata_60,afi_rdata_59,
afi_rdata_58,afi_rdata_57,afi_rdata_56,afi_rdata_55,afi_rdata_54,afi_rdata_53,afi_rdata_52,afi_rdata_51,afi_rdata_50,afi_rdata_49,afi_rdata_48,afi_rdata_47,afi_rdata_46,afi_rdata_45,afi_rdata_44,afi_rdata_43,afi_rdata_42,afi_rdata_41,afi_rdata_40,afi_rdata_39,afi_rdata_38,
afi_rdata_37,afi_rdata_36,afi_rdata_35,afi_rdata_34,afi_rdata_33,afi_rdata_32,afi_rdata_31,afi_rdata_30,afi_rdata_29,afi_rdata_28,afi_rdata_27,afi_rdata_26,afi_rdata_25,afi_rdata_24,afi_rdata_23,afi_rdata_22,afi_rdata_21,afi_rdata_20,afi_rdata_19,afi_rdata_18,afi_rdata_17,
afi_rdata_16,afi_rdata_15,afi_rdata_14,afi_rdata_13,afi_rdata_12,afi_rdata_11,afi_rdata_10,afi_rdata_9,afi_rdata_8,afi_rdata_7,afi_rdata_6,afi_rdata_5,afi_rdata_4,afi_rdata_3,afi_rdata_2,afi_rdata_1,afi_rdata_0}),
	.afi_wlat({afi_wlat_3,afi_wlat_2,afi_wlat_1,afi_wlat_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n({afi_cas_n_0}),
	.afi_ras_n({afi_ras_n_0}),
	.afi_rst_n({afi_rst_n_0}),
	.afi_we_n({afi_we_n_0}),
	.afi_addr({afi_addr_19,afi_addr_18,afi_addr_17,afi_addr_16,afi_addr_15,afi_addr_14,afi_addr_13,afi_addr_12,afi_addr_11,afi_addr_10,afi_addr_9,afi_addr_8,afi_addr_7,afi_addr_6,afi_addr_5,afi_addr_4,afi_addr_3,afi_addr_2,afi_addr_1,afi_addr_0}),
	.afi_ba({afi_ba_2,afi_ba_1,afi_ba_0}),
	.afi_cke({afi_cke_1,afi_cke_0}),
	.afi_cs_n({afi_cs_n_1,afi_cs_n_0}),
	.afi_dm({afi_dm_int_9,afi_dm_int_8,afi_dm_int_7,afi_dm_int_6,afi_dm_int_5,afi_dm_int_4,afi_dm_int_3,afi_dm_int_2,afi_dm_int_1,afi_dm_int_0}),
	.afi_dqs_burst({afi_dqs_burst_4,afi_dqs_burst_3,afi_dqs_burst_2,afi_dqs_burst_1,afi_dqs_burst_0}),
	.afi_odt({afi_odt_1,afi_odt_0}),
	.afi_rdata_en({afi_rdata_en_4,afi_rdata_en_3,afi_rdata_en_2,afi_rdata_en_1,afi_rdata_en_0}),
	.afi_rdata_en_full({afi_rdata_en_full_4,afi_rdata_en_full_3,afi_rdata_en_full_2,afi_rdata_en_full_1,afi_rdata_en_full_0}),
	.afi_wdata({afi_wdata_int_79,afi_wdata_int_78,afi_wdata_int_77,afi_wdata_int_76,afi_wdata_int_75,afi_wdata_int_74,afi_wdata_int_73,afi_wdata_int_72,afi_wdata_int_71,afi_wdata_int_70,afi_wdata_int_69,afi_wdata_int_68,afi_wdata_int_67,afi_wdata_int_66,afi_wdata_int_65,afi_wdata_int_64,
afi_wdata_int_63,afi_wdata_int_62,afi_wdata_int_61,afi_wdata_int_60,afi_wdata_int_59,afi_wdata_int_58,afi_wdata_int_57,afi_wdata_int_56,afi_wdata_int_55,afi_wdata_int_54,afi_wdata_int_53,afi_wdata_int_52,afi_wdata_int_51,afi_wdata_int_50,afi_wdata_int_49,afi_wdata_int_48,
afi_wdata_int_47,afi_wdata_int_46,afi_wdata_int_45,afi_wdata_int_44,afi_wdata_int_43,afi_wdata_int_42,afi_wdata_int_41,afi_wdata_int_40,afi_wdata_int_39,afi_wdata_int_38,afi_wdata_int_37,afi_wdata_int_36,afi_wdata_int_35,afi_wdata_int_34,afi_wdata_int_33,afi_wdata_int_32,
afi_wdata_int_31,afi_wdata_int_30,afi_wdata_int_29,afi_wdata_int_28,afi_wdata_int_27,afi_wdata_int_26,afi_wdata_int_25,afi_wdata_int_24,afi_wdata_int_23,afi_wdata_int_22,afi_wdata_int_21,afi_wdata_int_20,afi_wdata_int_19,afi_wdata_int_18,afi_wdata_int_17,afi_wdata_int_16,
afi_wdata_int_15,afi_wdata_int_14,afi_wdata_int_13,afi_wdata_int_12,afi_wdata_int_11,afi_wdata_int_10,afi_wdata_int_9,afi_wdata_int_8,afi_wdata_int_7,afi_wdata_int_6,afi_wdata_int_5,afi_wdata_int_4,afi_wdata_int_3,afi_wdata_int_2,afi_wdata_int_1,afi_wdata_int_0}),
	.afi_wdata_valid({afi_wdata_valid_4,afi_wdata_valid_3,afi_wdata_valid_2,afi_wdata_valid_1,afi_wdata_valid_0}),
	.cfg_addlat({gnd,gnd,gnd,cfg_addlat_wire_4,cfg_addlat_wire_3,cfg_addlat_wire_2,cfg_addlat_wire_1,cfg_addlat_wire_0}),
	.cfg_bankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth_wire_2,cfg_bankaddrwidth_wire_1,cfg_bankaddrwidth_wire_0}),
	.cfg_caswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat_wire_3,cfg_caswrlat_wire_2,cfg_caswrlat_wire_1,cfg_caswrlat_wire_0}),
	.cfg_coladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth_wire_4,cfg_coladdrwidth_wire_3,cfg_coladdrwidth_wire_2,cfg_coladdrwidth_wire_1,cfg_coladdrwidth_wire_0}),
	.cfg_csaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth_wire_2,cfg_csaddrwidth_wire_1,cfg_csaddrwidth_wire_0}),
	.cfg_devicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth_wire_3,cfg_devicewidth_wire_2,cfg_devicewidth_wire_1,cfg_devicewidth_wire_0}),
	.cfg_interfacewidth({cfg_interfacewidth_wire_7,cfg_interfacewidth_wire_6,cfg_interfacewidth_wire_5,cfg_interfacewidth_wire_4,cfg_interfacewidth_wire_3,cfg_interfacewidth_wire_2,cfg_interfacewidth_wire_1,cfg_interfacewidth_wire_0}),
	.cfg_rowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth_wire_4,cfg_rowaddrwidth_wire_3,cfg_rowaddrwidth_wire_2,cfg_rowaddrwidth_wire_1,cfg_rowaddrwidth_wire_0}),
	.cfg_tcl({gnd,gnd,gnd,cfg_tcl_wire_4,cfg_tcl_wire_3,cfg_tcl_wire_2,cfg_tcl_wire_1,cfg_tcl_wire_0}),
	.cfg_tmrd({gnd,gnd,gnd,gnd,cfg_tmrd_wire_3,cfg_tmrd_wire_2,cfg_tmrd_wire_1,cfg_tmrd_wire_0}),
	.cfg_trefi({gnd,gnd,gnd,cfg_trefi_wire_12,cfg_trefi_wire_11,cfg_trefi_wire_10,cfg_trefi_wire_9,cfg_trefi_wire_8,cfg_trefi_wire_7,cfg_trefi_wire_6,cfg_trefi_wire_5,cfg_trefi_wire_4,cfg_trefi_wire_3,cfg_trefi_wire_2,cfg_trefi_wire_1,cfg_trefi_wire_0}),
	.cfg_trfc({cfg_trfc_wire_7,cfg_trfc_wire_6,cfg_trfc_wire_5,cfg_trfc_wire_4,cfg_trfc_wire_3,cfg_trfc_wire_2,cfg_trfc_wire_1,cfg_trfc_wire_0}),
	.cfg_twr({gnd,gnd,gnd,gnd,cfg_twr_wire_3,cfg_twr_wire_2,cfg_twr_wire_1,cfg_twr_wire_0}),
	.afi_mem_clk_disable({afi_mem_clk_disable_0}),
	.cfg_dramconfig({gnd,gnd,gnd,cfg_dramconfig_wire_20,cfg_dramconfig_wire_19,cfg_dramconfig_wire_18,cfg_dramconfig_wire_17,cfg_dramconfig_wire_16,cfg_dramconfig_wire_15,cfg_dramconfig_wire_14,cfg_dramconfig_wire_13,cfg_dramconfig_wire_12,cfg_dramconfig_wire_11,cfg_dramconfig_wire_10,
cfg_dramconfig_wire_9,cfg_dramconfig_wire_8,cfg_dramconfig_wire_7,cfg_dramconfig_wire_6,cfg_dramconfig_wire_5,cfg_dramconfig_wire_4,cfg_dramconfig_wire_3,cfg_dramconfig_wire_2,cfg_dramconfig_wire_1,cfg_dramconfig_wire_0}),
	.leveled_dqs_clocks_0(leveled_dqs_clocks_0),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module soc_system_hps_sdram_p0_acv_hard_memphy (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	leveled_dqs_clocks_0,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	[0:0] afi_rdata_valid;
output 	ctl_reset_n;
output 	[79:0] afi_rdata;
output 	[3:0] afi_wlat;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	[0:0] afi_cas_n;
input 	[0:0] afi_ras_n;
input 	[0:0] afi_rst_n;
input 	[0:0] afi_we_n;
input 	[19:0] afi_addr;
input 	[2:0] afi_ba;
input 	[1:0] afi_cke;
input 	[1:0] afi_cs_n;
input 	[9:0] afi_dm;
input 	[4:0] afi_dqs_burst;
input 	[1:0] afi_odt;
input 	[4:0] afi_rdata_en;
input 	[4:0] afi_rdata_en_full;
input 	[79:0] afi_wdata;
input 	[4:0] afi_wdata_valid;
input 	[7:0] cfg_addlat;
input 	[7:0] cfg_bankaddrwidth;
input 	[7:0] cfg_caswrlat;
input 	[7:0] cfg_coladdrwidth;
input 	[7:0] cfg_csaddrwidth;
input 	[7:0] cfg_devicewidth;
input 	[7:0] cfg_interfacewidth;
input 	[7:0] cfg_rowaddrwidth;
input 	[7:0] cfg_tcl;
input 	[7:0] cfg_tmrd;
input 	[15:0] cfg_trefi;
input 	[7:0] cfg_trfc;
input 	[7:0] cfg_twr;
input 	[0:0] afi_mem_clk_disable;
input 	[23:0] cfg_dramconfig;
output 	leveled_dqs_clocks_0;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \memphy_ldc|leveled_hr_clocks[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \phy_ddio_address[0] ;
wire \phy_ddio_address[1] ;
wire \phy_ddio_address[2] ;
wire \phy_ddio_address[3] ;
wire \phy_ddio_address[4] ;
wire \phy_ddio_address[5] ;
wire \phy_ddio_address[6] ;
wire \phy_ddio_address[7] ;
wire \phy_ddio_address[8] ;
wire \phy_ddio_address[9] ;
wire \phy_ddio_address[10] ;
wire \phy_ddio_address[11] ;
wire \phy_ddio_address[12] ;
wire \phy_ddio_address[13] ;
wire \phy_ddio_address[14] ;
wire \phy_ddio_address[15] ;
wire \phy_ddio_address[16] ;
wire \phy_ddio_address[17] ;
wire \phy_ddio_address[18] ;
wire \phy_ddio_address[19] ;
wire \phy_ddio_address[20] ;
wire \phy_ddio_address[21] ;
wire \phy_ddio_address[22] ;
wire \phy_ddio_address[23] ;
wire \phy_ddio_address[24] ;
wire \phy_ddio_address[25] ;
wire \phy_ddio_address[26] ;
wire \phy_ddio_address[27] ;
wire \phy_ddio_address[28] ;
wire \phy_ddio_address[29] ;
wire \phy_ddio_address[30] ;
wire \phy_ddio_address[31] ;
wire \phy_ddio_address[32] ;
wire \phy_ddio_address[33] ;
wire \phy_ddio_address[34] ;
wire \phy_ddio_address[35] ;
wire \phy_ddio_address[36] ;
wire \phy_ddio_address[37] ;
wire \phy_ddio_address[38] ;
wire \phy_ddio_address[39] ;
wire \phy_ddio_address[40] ;
wire \phy_ddio_address[41] ;
wire \phy_ddio_address[42] ;
wire \phy_ddio_address[43] ;
wire \phy_ddio_address[44] ;
wire \phy_ddio_address[45] ;
wire \phy_ddio_address[46] ;
wire \phy_ddio_address[47] ;
wire \phy_ddio_address[48] ;
wire \phy_ddio_address[49] ;
wire \phy_ddio_address[50] ;
wire \phy_ddio_address[51] ;
wire \phy_ddio_address[52] ;
wire \phy_ddio_address[53] ;
wire \phy_ddio_address[54] ;
wire \phy_ddio_address[55] ;
wire \phy_ddio_address[56] ;
wire \phy_ddio_address[57] ;
wire \phy_ddio_address[58] ;
wire \phy_ddio_address[59] ;
wire \phy_ddio_bank[0] ;
wire \phy_ddio_bank[1] ;
wire \phy_ddio_bank[2] ;
wire \phy_ddio_bank[3] ;
wire \phy_ddio_bank[4] ;
wire \phy_ddio_bank[5] ;
wire \phy_ddio_bank[6] ;
wire \phy_ddio_bank[7] ;
wire \phy_ddio_bank[8] ;
wire \phy_ddio_bank[9] ;
wire \phy_ddio_bank[10] ;
wire \phy_ddio_bank[11] ;
wire \phy_ddio_cas_n[0] ;
wire \phy_ddio_cas_n[1] ;
wire \phy_ddio_cas_n[2] ;
wire \phy_ddio_cas_n[3] ;
wire \phy_ddio_ck[0] ;
wire \phy_ddio_ck[1] ;
wire \phy_ddio_cke[0] ;
wire \phy_ddio_cke[1] ;
wire \phy_ddio_cke[2] ;
wire \phy_ddio_cke[3] ;
wire \phy_ddio_cs_n[0] ;
wire \phy_ddio_cs_n[1] ;
wire \phy_ddio_cs_n[2] ;
wire \phy_ddio_cs_n[3] ;
wire \phy_ddio_dmdout[0] ;
wire \phy_ddio_dmdout[1] ;
wire \phy_ddio_dmdout[2] ;
wire \phy_ddio_dmdout[3] ;
wire \phy_ddio_dmdout[4] ;
wire \phy_ddio_dmdout[5] ;
wire \phy_ddio_dmdout[6] ;
wire \phy_ddio_dmdout[7] ;
wire \phy_ddio_dmdout[8] ;
wire \phy_ddio_dmdout[9] ;
wire \phy_ddio_dmdout[10] ;
wire \phy_ddio_dmdout[11] ;
wire \phy_ddio_dmdout[12] ;
wire \phy_ddio_dmdout[13] ;
wire \phy_ddio_dmdout[14] ;
wire \phy_ddio_dmdout[15] ;
wire \phy_ddio_dqdout[0] ;
wire \phy_ddio_dqdout[1] ;
wire \phy_ddio_dqdout[2] ;
wire \phy_ddio_dqdout[3] ;
wire \phy_ddio_dqdout[4] ;
wire \phy_ddio_dqdout[5] ;
wire \phy_ddio_dqdout[6] ;
wire \phy_ddio_dqdout[7] ;
wire \phy_ddio_dqdout[8] ;
wire \phy_ddio_dqdout[9] ;
wire \phy_ddio_dqdout[10] ;
wire \phy_ddio_dqdout[11] ;
wire \phy_ddio_dqdout[12] ;
wire \phy_ddio_dqdout[13] ;
wire \phy_ddio_dqdout[14] ;
wire \phy_ddio_dqdout[15] ;
wire \phy_ddio_dqdout[16] ;
wire \phy_ddio_dqdout[17] ;
wire \phy_ddio_dqdout[18] ;
wire \phy_ddio_dqdout[19] ;
wire \phy_ddio_dqdout[20] ;
wire \phy_ddio_dqdout[21] ;
wire \phy_ddio_dqdout[22] ;
wire \phy_ddio_dqdout[23] ;
wire \phy_ddio_dqdout[24] ;
wire \phy_ddio_dqdout[25] ;
wire \phy_ddio_dqdout[26] ;
wire \phy_ddio_dqdout[27] ;
wire \phy_ddio_dqdout[28] ;
wire \phy_ddio_dqdout[29] ;
wire \phy_ddio_dqdout[30] ;
wire \phy_ddio_dqdout[31] ;
wire \phy_ddio_dqdout[36] ;
wire \phy_ddio_dqdout[37] ;
wire \phy_ddio_dqdout[38] ;
wire \phy_ddio_dqdout[39] ;
wire \phy_ddio_dqdout[40] ;
wire \phy_ddio_dqdout[41] ;
wire \phy_ddio_dqdout[42] ;
wire \phy_ddio_dqdout[43] ;
wire \phy_ddio_dqdout[44] ;
wire \phy_ddio_dqdout[45] ;
wire \phy_ddio_dqdout[46] ;
wire \phy_ddio_dqdout[47] ;
wire \phy_ddio_dqdout[48] ;
wire \phy_ddio_dqdout[49] ;
wire \phy_ddio_dqdout[50] ;
wire \phy_ddio_dqdout[51] ;
wire \phy_ddio_dqdout[52] ;
wire \phy_ddio_dqdout[53] ;
wire \phy_ddio_dqdout[54] ;
wire \phy_ddio_dqdout[55] ;
wire \phy_ddio_dqdout[56] ;
wire \phy_ddio_dqdout[57] ;
wire \phy_ddio_dqdout[58] ;
wire \phy_ddio_dqdout[59] ;
wire \phy_ddio_dqdout[60] ;
wire \phy_ddio_dqdout[61] ;
wire \phy_ddio_dqdout[62] ;
wire \phy_ddio_dqdout[63] ;
wire \phy_ddio_dqdout[64] ;
wire \phy_ddio_dqdout[65] ;
wire \phy_ddio_dqdout[66] ;
wire \phy_ddio_dqdout[67] ;
wire \phy_ddio_dqdout[72] ;
wire \phy_ddio_dqdout[73] ;
wire \phy_ddio_dqdout[74] ;
wire \phy_ddio_dqdout[75] ;
wire \phy_ddio_dqdout[76] ;
wire \phy_ddio_dqdout[77] ;
wire \phy_ddio_dqdout[78] ;
wire \phy_ddio_dqdout[79] ;
wire \phy_ddio_dqdout[80] ;
wire \phy_ddio_dqdout[81] ;
wire \phy_ddio_dqdout[82] ;
wire \phy_ddio_dqdout[83] ;
wire \phy_ddio_dqdout[84] ;
wire \phy_ddio_dqdout[85] ;
wire \phy_ddio_dqdout[86] ;
wire \phy_ddio_dqdout[87] ;
wire \phy_ddio_dqdout[88] ;
wire \phy_ddio_dqdout[89] ;
wire \phy_ddio_dqdout[90] ;
wire \phy_ddio_dqdout[91] ;
wire \phy_ddio_dqdout[92] ;
wire \phy_ddio_dqdout[93] ;
wire \phy_ddio_dqdout[94] ;
wire \phy_ddio_dqdout[95] ;
wire \phy_ddio_dqdout[96] ;
wire \phy_ddio_dqdout[97] ;
wire \phy_ddio_dqdout[98] ;
wire \phy_ddio_dqdout[99] ;
wire \phy_ddio_dqdout[100] ;
wire \phy_ddio_dqdout[101] ;
wire \phy_ddio_dqdout[102] ;
wire \phy_ddio_dqdout[103] ;
wire \phy_ddio_dqdout[108] ;
wire \phy_ddio_dqdout[109] ;
wire \phy_ddio_dqdout[110] ;
wire \phy_ddio_dqdout[111] ;
wire \phy_ddio_dqdout[112] ;
wire \phy_ddio_dqdout[113] ;
wire \phy_ddio_dqdout[114] ;
wire \phy_ddio_dqdout[115] ;
wire \phy_ddio_dqdout[116] ;
wire \phy_ddio_dqdout[117] ;
wire \phy_ddio_dqdout[118] ;
wire \phy_ddio_dqdout[119] ;
wire \phy_ddio_dqdout[120] ;
wire \phy_ddio_dqdout[121] ;
wire \phy_ddio_dqdout[122] ;
wire \phy_ddio_dqdout[123] ;
wire \phy_ddio_dqdout[124] ;
wire \phy_ddio_dqdout[125] ;
wire \phy_ddio_dqdout[126] ;
wire \phy_ddio_dqdout[127] ;
wire \phy_ddio_dqdout[128] ;
wire \phy_ddio_dqdout[129] ;
wire \phy_ddio_dqdout[130] ;
wire \phy_ddio_dqdout[131] ;
wire \phy_ddio_dqdout[132] ;
wire \phy_ddio_dqdout[133] ;
wire \phy_ddio_dqdout[134] ;
wire \phy_ddio_dqdout[135] ;
wire \phy_ddio_dqdout[136] ;
wire \phy_ddio_dqdout[137] ;
wire \phy_ddio_dqdout[138] ;
wire \phy_ddio_dqdout[139] ;
wire \phy_ddio_dqoe[0] ;
wire \phy_ddio_dqoe[1] ;
wire \phy_ddio_dqoe[2] ;
wire \phy_ddio_dqoe[3] ;
wire \phy_ddio_dqoe[4] ;
wire \phy_ddio_dqoe[5] ;
wire \phy_ddio_dqoe[6] ;
wire \phy_ddio_dqoe[7] ;
wire \phy_ddio_dqoe[8] ;
wire \phy_ddio_dqoe[9] ;
wire \phy_ddio_dqoe[10] ;
wire \phy_ddio_dqoe[11] ;
wire \phy_ddio_dqoe[12] ;
wire \phy_ddio_dqoe[13] ;
wire \phy_ddio_dqoe[14] ;
wire \phy_ddio_dqoe[15] ;
wire \phy_ddio_dqoe[18] ;
wire \phy_ddio_dqoe[19] ;
wire \phy_ddio_dqoe[20] ;
wire \phy_ddio_dqoe[21] ;
wire \phy_ddio_dqoe[22] ;
wire \phy_ddio_dqoe[23] ;
wire \phy_ddio_dqoe[24] ;
wire \phy_ddio_dqoe[25] ;
wire \phy_ddio_dqoe[26] ;
wire \phy_ddio_dqoe[27] ;
wire \phy_ddio_dqoe[28] ;
wire \phy_ddio_dqoe[29] ;
wire \phy_ddio_dqoe[30] ;
wire \phy_ddio_dqoe[31] ;
wire \phy_ddio_dqoe[32] ;
wire \phy_ddio_dqoe[33] ;
wire \phy_ddio_dqoe[36] ;
wire \phy_ddio_dqoe[37] ;
wire \phy_ddio_dqoe[38] ;
wire \phy_ddio_dqoe[39] ;
wire \phy_ddio_dqoe[40] ;
wire \phy_ddio_dqoe[41] ;
wire \phy_ddio_dqoe[42] ;
wire \phy_ddio_dqoe[43] ;
wire \phy_ddio_dqoe[44] ;
wire \phy_ddio_dqoe[45] ;
wire \phy_ddio_dqoe[46] ;
wire \phy_ddio_dqoe[47] ;
wire \phy_ddio_dqoe[48] ;
wire \phy_ddio_dqoe[49] ;
wire \phy_ddio_dqoe[50] ;
wire \phy_ddio_dqoe[51] ;
wire \phy_ddio_dqoe[54] ;
wire \phy_ddio_dqoe[55] ;
wire \phy_ddio_dqoe[56] ;
wire \phy_ddio_dqoe[57] ;
wire \phy_ddio_dqoe[58] ;
wire \phy_ddio_dqoe[59] ;
wire \phy_ddio_dqoe[60] ;
wire \phy_ddio_dqoe[61] ;
wire \phy_ddio_dqoe[62] ;
wire \phy_ddio_dqoe[63] ;
wire \phy_ddio_dqoe[64] ;
wire \phy_ddio_dqoe[65] ;
wire \phy_ddio_dqoe[66] ;
wire \phy_ddio_dqoe[67] ;
wire \phy_ddio_dqoe[68] ;
wire \phy_ddio_dqoe[69] ;
wire \phy_ddio_dqs_dout[0] ;
wire \phy_ddio_dqs_dout[1] ;
wire \phy_ddio_dqs_dout[2] ;
wire \phy_ddio_dqs_dout[3] ;
wire \phy_ddio_dqs_dout[4] ;
wire \phy_ddio_dqs_dout[5] ;
wire \phy_ddio_dqs_dout[6] ;
wire \phy_ddio_dqs_dout[7] ;
wire \phy_ddio_dqs_dout[8] ;
wire \phy_ddio_dqs_dout[9] ;
wire \phy_ddio_dqs_dout[10] ;
wire \phy_ddio_dqs_dout[11] ;
wire \phy_ddio_dqs_dout[12] ;
wire \phy_ddio_dqs_dout[13] ;
wire \phy_ddio_dqs_dout[14] ;
wire \phy_ddio_dqs_dout[15] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[0] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[1] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[2] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[3] ;
wire \phy_ddio_dqslogic_aclr_pstamble[0] ;
wire \phy_ddio_dqslogic_aclr_pstamble[1] ;
wire \phy_ddio_dqslogic_aclr_pstamble[2] ;
wire \phy_ddio_dqslogic_aclr_pstamble[3] ;
wire \phy_ddio_dqslogic_dqsena[0] ;
wire \phy_ddio_dqslogic_dqsena[1] ;
wire \phy_ddio_dqslogic_dqsena[2] ;
wire \phy_ddio_dqslogic_dqsena[3] ;
wire \phy_ddio_dqslogic_dqsena[4] ;
wire \phy_ddio_dqslogic_dqsena[5] ;
wire \phy_ddio_dqslogic_dqsena[6] ;
wire \phy_ddio_dqslogic_dqsena[7] ;
wire \phy_ddio_dqslogic_fiforeset[0] ;
wire \phy_ddio_dqslogic_fiforeset[1] ;
wire \phy_ddio_dqslogic_fiforeset[2] ;
wire \phy_ddio_dqslogic_fiforeset[3] ;
wire \phy_ddio_dqslogic_incrdataen[0] ;
wire \phy_ddio_dqslogic_incrdataen[1] ;
wire \phy_ddio_dqslogic_incrdataen[2] ;
wire \phy_ddio_dqslogic_incrdataen[3] ;
wire \phy_ddio_dqslogic_incrdataen[4] ;
wire \phy_ddio_dqslogic_incrdataen[5] ;
wire \phy_ddio_dqslogic_incrdataen[6] ;
wire \phy_ddio_dqslogic_incrdataen[7] ;
wire \phy_ddio_dqslogic_incwrptr[0] ;
wire \phy_ddio_dqslogic_incwrptr[1] ;
wire \phy_ddio_dqslogic_incwrptr[2] ;
wire \phy_ddio_dqslogic_incwrptr[3] ;
wire \phy_ddio_dqslogic_incwrptr[4] ;
wire \phy_ddio_dqslogic_incwrptr[5] ;
wire \phy_ddio_dqslogic_incwrptr[6] ;
wire \phy_ddio_dqslogic_incwrptr[7] ;
wire \phy_ddio_dqslogic_oct[0] ;
wire \phy_ddio_dqslogic_oct[1] ;
wire \phy_ddio_dqslogic_oct[2] ;
wire \phy_ddio_dqslogic_oct[3] ;
wire \phy_ddio_dqslogic_oct[4] ;
wire \phy_ddio_dqslogic_oct[5] ;
wire \phy_ddio_dqslogic_oct[6] ;
wire \phy_ddio_dqslogic_oct[7] ;
wire \phy_ddio_dqslogic_readlatency[0] ;
wire \phy_ddio_dqslogic_readlatency[1] ;
wire \phy_ddio_dqslogic_readlatency[2] ;
wire \phy_ddio_dqslogic_readlatency[3] ;
wire \phy_ddio_dqslogic_readlatency[4] ;
wire \phy_ddio_dqslogic_readlatency[5] ;
wire \phy_ddio_dqslogic_readlatency[6] ;
wire \phy_ddio_dqslogic_readlatency[7] ;
wire \phy_ddio_dqslogic_readlatency[8] ;
wire \phy_ddio_dqslogic_readlatency[9] ;
wire \phy_ddio_dqslogic_readlatency[10] ;
wire \phy_ddio_dqslogic_readlatency[11] ;
wire \phy_ddio_dqslogic_readlatency[12] ;
wire \phy_ddio_dqslogic_readlatency[13] ;
wire \phy_ddio_dqslogic_readlatency[14] ;
wire \phy_ddio_dqslogic_readlatency[15] ;
wire \phy_ddio_dqslogic_readlatency[16] ;
wire \phy_ddio_dqslogic_readlatency[17] ;
wire \phy_ddio_dqslogic_readlatency[18] ;
wire \phy_ddio_dqslogic_readlatency[19] ;
wire \phy_ddio_dqs_oe[0] ;
wire \phy_ddio_dqs_oe[1] ;
wire \phy_ddio_dqs_oe[2] ;
wire \phy_ddio_dqs_oe[3] ;
wire \phy_ddio_dqs_oe[4] ;
wire \phy_ddio_dqs_oe[5] ;
wire \phy_ddio_dqs_oe[6] ;
wire \phy_ddio_dqs_oe[7] ;
wire \phy_ddio_odt[0] ;
wire \phy_ddio_odt[1] ;
wire \phy_ddio_odt[2] ;
wire \phy_ddio_odt[3] ;
wire \phy_ddio_ras_n[0] ;
wire \phy_ddio_ras_n[1] ;
wire \phy_ddio_ras_n[2] ;
wire \phy_ddio_ras_n[3] ;
wire \phy_ddio_reset_n[0] ;
wire \phy_ddio_reset_n[1] ;
wire \phy_ddio_reset_n[2] ;
wire \phy_ddio_reset_n[3] ;
wire \phy_ddio_we_n[0] ;
wire \phy_ddio_we_n[1] ;
wire \phy_ddio_we_n[2] ;
wire \phy_ddio_we_n[3] ;

wire [79:0] hphy_inst_AFIRDATA_bus;
wire [3:0] hphy_inst_AFIWLAT_bus;
wire [63:0] hphy_inst_PHYDDIOADDRDOUT_bus;
wire [11:0] hphy_inst_PHYDDIOBADOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCKDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCKEDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCSNDOUT_bus;
wire [19:0] hphy_inst_PHYDDIODMDOUT_bus;
wire [179:0] hphy_inst_PHYDDIODQDOUT_bus;
wire [89:0] hphy_inst_PHYDDIODQOE_bus;
wire [19:0] hphy_inst_PHYDDIODQSDOUT_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICDQSENA_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICFIFORESET_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICOCT_bus;
wire [24:0] hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus;
wire [9:0] hphy_inst_PHYDDIODQSOE_bus;
wire [7:0] hphy_inst_PHYDDIOODTDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORESETNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOWENDOUT_bus;

assign afi_rdata[0] = hphy_inst_AFIRDATA_bus[0];
assign afi_rdata[1] = hphy_inst_AFIRDATA_bus[1];
assign afi_rdata[2] = hphy_inst_AFIRDATA_bus[2];
assign afi_rdata[3] = hphy_inst_AFIRDATA_bus[3];
assign afi_rdata[4] = hphy_inst_AFIRDATA_bus[4];
assign afi_rdata[5] = hphy_inst_AFIRDATA_bus[5];
assign afi_rdata[6] = hphy_inst_AFIRDATA_bus[6];
assign afi_rdata[7] = hphy_inst_AFIRDATA_bus[7];
assign afi_rdata[8] = hphy_inst_AFIRDATA_bus[8];
assign afi_rdata[9] = hphy_inst_AFIRDATA_bus[9];
assign afi_rdata[10] = hphy_inst_AFIRDATA_bus[10];
assign afi_rdata[11] = hphy_inst_AFIRDATA_bus[11];
assign afi_rdata[12] = hphy_inst_AFIRDATA_bus[12];
assign afi_rdata[13] = hphy_inst_AFIRDATA_bus[13];
assign afi_rdata[14] = hphy_inst_AFIRDATA_bus[14];
assign afi_rdata[15] = hphy_inst_AFIRDATA_bus[15];
assign afi_rdata[16] = hphy_inst_AFIRDATA_bus[16];
assign afi_rdata[17] = hphy_inst_AFIRDATA_bus[17];
assign afi_rdata[18] = hphy_inst_AFIRDATA_bus[18];
assign afi_rdata[19] = hphy_inst_AFIRDATA_bus[19];
assign afi_rdata[20] = hphy_inst_AFIRDATA_bus[20];
assign afi_rdata[21] = hphy_inst_AFIRDATA_bus[21];
assign afi_rdata[22] = hphy_inst_AFIRDATA_bus[22];
assign afi_rdata[23] = hphy_inst_AFIRDATA_bus[23];
assign afi_rdata[24] = hphy_inst_AFIRDATA_bus[24];
assign afi_rdata[25] = hphy_inst_AFIRDATA_bus[25];
assign afi_rdata[26] = hphy_inst_AFIRDATA_bus[26];
assign afi_rdata[27] = hphy_inst_AFIRDATA_bus[27];
assign afi_rdata[28] = hphy_inst_AFIRDATA_bus[28];
assign afi_rdata[29] = hphy_inst_AFIRDATA_bus[29];
assign afi_rdata[30] = hphy_inst_AFIRDATA_bus[30];
assign afi_rdata[31] = hphy_inst_AFIRDATA_bus[31];
assign afi_rdata[32] = hphy_inst_AFIRDATA_bus[32];
assign afi_rdata[33] = hphy_inst_AFIRDATA_bus[33];
assign afi_rdata[34] = hphy_inst_AFIRDATA_bus[34];
assign afi_rdata[35] = hphy_inst_AFIRDATA_bus[35];
assign afi_rdata[36] = hphy_inst_AFIRDATA_bus[36];
assign afi_rdata[37] = hphy_inst_AFIRDATA_bus[37];
assign afi_rdata[38] = hphy_inst_AFIRDATA_bus[38];
assign afi_rdata[39] = hphy_inst_AFIRDATA_bus[39];
assign afi_rdata[40] = hphy_inst_AFIRDATA_bus[40];
assign afi_rdata[41] = hphy_inst_AFIRDATA_bus[41];
assign afi_rdata[42] = hphy_inst_AFIRDATA_bus[42];
assign afi_rdata[43] = hphy_inst_AFIRDATA_bus[43];
assign afi_rdata[44] = hphy_inst_AFIRDATA_bus[44];
assign afi_rdata[45] = hphy_inst_AFIRDATA_bus[45];
assign afi_rdata[46] = hphy_inst_AFIRDATA_bus[46];
assign afi_rdata[47] = hphy_inst_AFIRDATA_bus[47];
assign afi_rdata[48] = hphy_inst_AFIRDATA_bus[48];
assign afi_rdata[49] = hphy_inst_AFIRDATA_bus[49];
assign afi_rdata[50] = hphy_inst_AFIRDATA_bus[50];
assign afi_rdata[51] = hphy_inst_AFIRDATA_bus[51];
assign afi_rdata[52] = hphy_inst_AFIRDATA_bus[52];
assign afi_rdata[53] = hphy_inst_AFIRDATA_bus[53];
assign afi_rdata[54] = hphy_inst_AFIRDATA_bus[54];
assign afi_rdata[55] = hphy_inst_AFIRDATA_bus[55];
assign afi_rdata[56] = hphy_inst_AFIRDATA_bus[56];
assign afi_rdata[57] = hphy_inst_AFIRDATA_bus[57];
assign afi_rdata[58] = hphy_inst_AFIRDATA_bus[58];
assign afi_rdata[59] = hphy_inst_AFIRDATA_bus[59];
assign afi_rdata[60] = hphy_inst_AFIRDATA_bus[60];
assign afi_rdata[61] = hphy_inst_AFIRDATA_bus[61];
assign afi_rdata[62] = hphy_inst_AFIRDATA_bus[62];
assign afi_rdata[63] = hphy_inst_AFIRDATA_bus[63];
assign afi_rdata[64] = hphy_inst_AFIRDATA_bus[64];
assign afi_rdata[65] = hphy_inst_AFIRDATA_bus[65];
assign afi_rdata[66] = hphy_inst_AFIRDATA_bus[66];
assign afi_rdata[67] = hphy_inst_AFIRDATA_bus[67];
assign afi_rdata[68] = hphy_inst_AFIRDATA_bus[68];
assign afi_rdata[69] = hphy_inst_AFIRDATA_bus[69];
assign afi_rdata[70] = hphy_inst_AFIRDATA_bus[70];
assign afi_rdata[71] = hphy_inst_AFIRDATA_bus[71];
assign afi_rdata[72] = hphy_inst_AFIRDATA_bus[72];
assign afi_rdata[73] = hphy_inst_AFIRDATA_bus[73];
assign afi_rdata[74] = hphy_inst_AFIRDATA_bus[74];
assign afi_rdata[75] = hphy_inst_AFIRDATA_bus[75];
assign afi_rdata[76] = hphy_inst_AFIRDATA_bus[76];
assign afi_rdata[77] = hphy_inst_AFIRDATA_bus[77];
assign afi_rdata[78] = hphy_inst_AFIRDATA_bus[78];
assign afi_rdata[79] = hphy_inst_AFIRDATA_bus[79];

assign afi_wlat[0] = hphy_inst_AFIWLAT_bus[0];
assign afi_wlat[1] = hphy_inst_AFIWLAT_bus[1];
assign afi_wlat[2] = hphy_inst_AFIWLAT_bus[2];
assign afi_wlat[3] = hphy_inst_AFIWLAT_bus[3];

assign \phy_ddio_address[0]  = hphy_inst_PHYDDIOADDRDOUT_bus[0];
assign \phy_ddio_address[1]  = hphy_inst_PHYDDIOADDRDOUT_bus[1];
assign \phy_ddio_address[2]  = hphy_inst_PHYDDIOADDRDOUT_bus[2];
assign \phy_ddio_address[3]  = hphy_inst_PHYDDIOADDRDOUT_bus[3];
assign \phy_ddio_address[4]  = hphy_inst_PHYDDIOADDRDOUT_bus[4];
assign \phy_ddio_address[5]  = hphy_inst_PHYDDIOADDRDOUT_bus[5];
assign \phy_ddio_address[6]  = hphy_inst_PHYDDIOADDRDOUT_bus[6];
assign \phy_ddio_address[7]  = hphy_inst_PHYDDIOADDRDOUT_bus[7];
assign \phy_ddio_address[8]  = hphy_inst_PHYDDIOADDRDOUT_bus[8];
assign \phy_ddio_address[9]  = hphy_inst_PHYDDIOADDRDOUT_bus[9];
assign \phy_ddio_address[10]  = hphy_inst_PHYDDIOADDRDOUT_bus[10];
assign \phy_ddio_address[11]  = hphy_inst_PHYDDIOADDRDOUT_bus[11];
assign \phy_ddio_address[12]  = hphy_inst_PHYDDIOADDRDOUT_bus[12];
assign \phy_ddio_address[13]  = hphy_inst_PHYDDIOADDRDOUT_bus[13];
assign \phy_ddio_address[14]  = hphy_inst_PHYDDIOADDRDOUT_bus[14];
assign \phy_ddio_address[15]  = hphy_inst_PHYDDIOADDRDOUT_bus[15];
assign \phy_ddio_address[16]  = hphy_inst_PHYDDIOADDRDOUT_bus[16];
assign \phy_ddio_address[17]  = hphy_inst_PHYDDIOADDRDOUT_bus[17];
assign \phy_ddio_address[18]  = hphy_inst_PHYDDIOADDRDOUT_bus[18];
assign \phy_ddio_address[19]  = hphy_inst_PHYDDIOADDRDOUT_bus[19];
assign \phy_ddio_address[20]  = hphy_inst_PHYDDIOADDRDOUT_bus[20];
assign \phy_ddio_address[21]  = hphy_inst_PHYDDIOADDRDOUT_bus[21];
assign \phy_ddio_address[22]  = hphy_inst_PHYDDIOADDRDOUT_bus[22];
assign \phy_ddio_address[23]  = hphy_inst_PHYDDIOADDRDOUT_bus[23];
assign \phy_ddio_address[24]  = hphy_inst_PHYDDIOADDRDOUT_bus[24];
assign \phy_ddio_address[25]  = hphy_inst_PHYDDIOADDRDOUT_bus[25];
assign \phy_ddio_address[26]  = hphy_inst_PHYDDIOADDRDOUT_bus[26];
assign \phy_ddio_address[27]  = hphy_inst_PHYDDIOADDRDOUT_bus[27];
assign \phy_ddio_address[28]  = hphy_inst_PHYDDIOADDRDOUT_bus[28];
assign \phy_ddio_address[29]  = hphy_inst_PHYDDIOADDRDOUT_bus[29];
assign \phy_ddio_address[30]  = hphy_inst_PHYDDIOADDRDOUT_bus[30];
assign \phy_ddio_address[31]  = hphy_inst_PHYDDIOADDRDOUT_bus[31];
assign \phy_ddio_address[32]  = hphy_inst_PHYDDIOADDRDOUT_bus[32];
assign \phy_ddio_address[33]  = hphy_inst_PHYDDIOADDRDOUT_bus[33];
assign \phy_ddio_address[34]  = hphy_inst_PHYDDIOADDRDOUT_bus[34];
assign \phy_ddio_address[35]  = hphy_inst_PHYDDIOADDRDOUT_bus[35];
assign \phy_ddio_address[36]  = hphy_inst_PHYDDIOADDRDOUT_bus[36];
assign \phy_ddio_address[37]  = hphy_inst_PHYDDIOADDRDOUT_bus[37];
assign \phy_ddio_address[38]  = hphy_inst_PHYDDIOADDRDOUT_bus[38];
assign \phy_ddio_address[39]  = hphy_inst_PHYDDIOADDRDOUT_bus[39];
assign \phy_ddio_address[40]  = hphy_inst_PHYDDIOADDRDOUT_bus[40];
assign \phy_ddio_address[41]  = hphy_inst_PHYDDIOADDRDOUT_bus[41];
assign \phy_ddio_address[42]  = hphy_inst_PHYDDIOADDRDOUT_bus[42];
assign \phy_ddio_address[43]  = hphy_inst_PHYDDIOADDRDOUT_bus[43];
assign \phy_ddio_address[44]  = hphy_inst_PHYDDIOADDRDOUT_bus[44];
assign \phy_ddio_address[45]  = hphy_inst_PHYDDIOADDRDOUT_bus[45];
assign \phy_ddio_address[46]  = hphy_inst_PHYDDIOADDRDOUT_bus[46];
assign \phy_ddio_address[47]  = hphy_inst_PHYDDIOADDRDOUT_bus[47];
assign \phy_ddio_address[48]  = hphy_inst_PHYDDIOADDRDOUT_bus[48];
assign \phy_ddio_address[49]  = hphy_inst_PHYDDIOADDRDOUT_bus[49];
assign \phy_ddio_address[50]  = hphy_inst_PHYDDIOADDRDOUT_bus[50];
assign \phy_ddio_address[51]  = hphy_inst_PHYDDIOADDRDOUT_bus[51];
assign \phy_ddio_address[52]  = hphy_inst_PHYDDIOADDRDOUT_bus[52];
assign \phy_ddio_address[53]  = hphy_inst_PHYDDIOADDRDOUT_bus[53];
assign \phy_ddio_address[54]  = hphy_inst_PHYDDIOADDRDOUT_bus[54];
assign \phy_ddio_address[55]  = hphy_inst_PHYDDIOADDRDOUT_bus[55];
assign \phy_ddio_address[56]  = hphy_inst_PHYDDIOADDRDOUT_bus[56];
assign \phy_ddio_address[57]  = hphy_inst_PHYDDIOADDRDOUT_bus[57];
assign \phy_ddio_address[58]  = hphy_inst_PHYDDIOADDRDOUT_bus[58];
assign \phy_ddio_address[59]  = hphy_inst_PHYDDIOADDRDOUT_bus[59];

assign \phy_ddio_bank[0]  = hphy_inst_PHYDDIOBADOUT_bus[0];
assign \phy_ddio_bank[1]  = hphy_inst_PHYDDIOBADOUT_bus[1];
assign \phy_ddio_bank[2]  = hphy_inst_PHYDDIOBADOUT_bus[2];
assign \phy_ddio_bank[3]  = hphy_inst_PHYDDIOBADOUT_bus[3];
assign \phy_ddio_bank[4]  = hphy_inst_PHYDDIOBADOUT_bus[4];
assign \phy_ddio_bank[5]  = hphy_inst_PHYDDIOBADOUT_bus[5];
assign \phy_ddio_bank[6]  = hphy_inst_PHYDDIOBADOUT_bus[6];
assign \phy_ddio_bank[7]  = hphy_inst_PHYDDIOBADOUT_bus[7];
assign \phy_ddio_bank[8]  = hphy_inst_PHYDDIOBADOUT_bus[8];
assign \phy_ddio_bank[9]  = hphy_inst_PHYDDIOBADOUT_bus[9];
assign \phy_ddio_bank[10]  = hphy_inst_PHYDDIOBADOUT_bus[10];
assign \phy_ddio_bank[11]  = hphy_inst_PHYDDIOBADOUT_bus[11];

assign \phy_ddio_cas_n[0]  = hphy_inst_PHYDDIOCASNDOUT_bus[0];
assign \phy_ddio_cas_n[1]  = hphy_inst_PHYDDIOCASNDOUT_bus[1];
assign \phy_ddio_cas_n[2]  = hphy_inst_PHYDDIOCASNDOUT_bus[2];
assign \phy_ddio_cas_n[3]  = hphy_inst_PHYDDIOCASNDOUT_bus[3];

assign \phy_ddio_ck[0]  = hphy_inst_PHYDDIOCKDOUT_bus[0];
assign \phy_ddio_ck[1]  = hphy_inst_PHYDDIOCKDOUT_bus[1];

assign \phy_ddio_cke[0]  = hphy_inst_PHYDDIOCKEDOUT_bus[0];
assign \phy_ddio_cke[1]  = hphy_inst_PHYDDIOCKEDOUT_bus[1];
assign \phy_ddio_cke[2]  = hphy_inst_PHYDDIOCKEDOUT_bus[2];
assign \phy_ddio_cke[3]  = hphy_inst_PHYDDIOCKEDOUT_bus[3];

assign \phy_ddio_cs_n[0]  = hphy_inst_PHYDDIOCSNDOUT_bus[0];
assign \phy_ddio_cs_n[1]  = hphy_inst_PHYDDIOCSNDOUT_bus[1];
assign \phy_ddio_cs_n[2]  = hphy_inst_PHYDDIOCSNDOUT_bus[2];
assign \phy_ddio_cs_n[3]  = hphy_inst_PHYDDIOCSNDOUT_bus[3];

assign \phy_ddio_dmdout[0]  = hphy_inst_PHYDDIODMDOUT_bus[0];
assign \phy_ddio_dmdout[1]  = hphy_inst_PHYDDIODMDOUT_bus[1];
assign \phy_ddio_dmdout[2]  = hphy_inst_PHYDDIODMDOUT_bus[2];
assign \phy_ddio_dmdout[3]  = hphy_inst_PHYDDIODMDOUT_bus[3];
assign \phy_ddio_dmdout[4]  = hphy_inst_PHYDDIODMDOUT_bus[4];
assign \phy_ddio_dmdout[5]  = hphy_inst_PHYDDIODMDOUT_bus[5];
assign \phy_ddio_dmdout[6]  = hphy_inst_PHYDDIODMDOUT_bus[6];
assign \phy_ddio_dmdout[7]  = hphy_inst_PHYDDIODMDOUT_bus[7];
assign \phy_ddio_dmdout[8]  = hphy_inst_PHYDDIODMDOUT_bus[8];
assign \phy_ddio_dmdout[9]  = hphy_inst_PHYDDIODMDOUT_bus[9];
assign \phy_ddio_dmdout[10]  = hphy_inst_PHYDDIODMDOUT_bus[10];
assign \phy_ddio_dmdout[11]  = hphy_inst_PHYDDIODMDOUT_bus[11];
assign \phy_ddio_dmdout[12]  = hphy_inst_PHYDDIODMDOUT_bus[12];
assign \phy_ddio_dmdout[13]  = hphy_inst_PHYDDIODMDOUT_bus[13];
assign \phy_ddio_dmdout[14]  = hphy_inst_PHYDDIODMDOUT_bus[14];
assign \phy_ddio_dmdout[15]  = hphy_inst_PHYDDIODMDOUT_bus[15];

assign \phy_ddio_dqdout[0]  = hphy_inst_PHYDDIODQDOUT_bus[0];
assign \phy_ddio_dqdout[1]  = hphy_inst_PHYDDIODQDOUT_bus[1];
assign \phy_ddio_dqdout[2]  = hphy_inst_PHYDDIODQDOUT_bus[2];
assign \phy_ddio_dqdout[3]  = hphy_inst_PHYDDIODQDOUT_bus[3];
assign \phy_ddio_dqdout[4]  = hphy_inst_PHYDDIODQDOUT_bus[4];
assign \phy_ddio_dqdout[5]  = hphy_inst_PHYDDIODQDOUT_bus[5];
assign \phy_ddio_dqdout[6]  = hphy_inst_PHYDDIODQDOUT_bus[6];
assign \phy_ddio_dqdout[7]  = hphy_inst_PHYDDIODQDOUT_bus[7];
assign \phy_ddio_dqdout[8]  = hphy_inst_PHYDDIODQDOUT_bus[8];
assign \phy_ddio_dqdout[9]  = hphy_inst_PHYDDIODQDOUT_bus[9];
assign \phy_ddio_dqdout[10]  = hphy_inst_PHYDDIODQDOUT_bus[10];
assign \phy_ddio_dqdout[11]  = hphy_inst_PHYDDIODQDOUT_bus[11];
assign \phy_ddio_dqdout[12]  = hphy_inst_PHYDDIODQDOUT_bus[12];
assign \phy_ddio_dqdout[13]  = hphy_inst_PHYDDIODQDOUT_bus[13];
assign \phy_ddio_dqdout[14]  = hphy_inst_PHYDDIODQDOUT_bus[14];
assign \phy_ddio_dqdout[15]  = hphy_inst_PHYDDIODQDOUT_bus[15];
assign \phy_ddio_dqdout[16]  = hphy_inst_PHYDDIODQDOUT_bus[16];
assign \phy_ddio_dqdout[17]  = hphy_inst_PHYDDIODQDOUT_bus[17];
assign \phy_ddio_dqdout[18]  = hphy_inst_PHYDDIODQDOUT_bus[18];
assign \phy_ddio_dqdout[19]  = hphy_inst_PHYDDIODQDOUT_bus[19];
assign \phy_ddio_dqdout[20]  = hphy_inst_PHYDDIODQDOUT_bus[20];
assign \phy_ddio_dqdout[21]  = hphy_inst_PHYDDIODQDOUT_bus[21];
assign \phy_ddio_dqdout[22]  = hphy_inst_PHYDDIODQDOUT_bus[22];
assign \phy_ddio_dqdout[23]  = hphy_inst_PHYDDIODQDOUT_bus[23];
assign \phy_ddio_dqdout[24]  = hphy_inst_PHYDDIODQDOUT_bus[24];
assign \phy_ddio_dqdout[25]  = hphy_inst_PHYDDIODQDOUT_bus[25];
assign \phy_ddio_dqdout[26]  = hphy_inst_PHYDDIODQDOUT_bus[26];
assign \phy_ddio_dqdout[27]  = hphy_inst_PHYDDIODQDOUT_bus[27];
assign \phy_ddio_dqdout[28]  = hphy_inst_PHYDDIODQDOUT_bus[28];
assign \phy_ddio_dqdout[29]  = hphy_inst_PHYDDIODQDOUT_bus[29];
assign \phy_ddio_dqdout[30]  = hphy_inst_PHYDDIODQDOUT_bus[30];
assign \phy_ddio_dqdout[31]  = hphy_inst_PHYDDIODQDOUT_bus[31];
assign \phy_ddio_dqdout[36]  = hphy_inst_PHYDDIODQDOUT_bus[36];
assign \phy_ddio_dqdout[37]  = hphy_inst_PHYDDIODQDOUT_bus[37];
assign \phy_ddio_dqdout[38]  = hphy_inst_PHYDDIODQDOUT_bus[38];
assign \phy_ddio_dqdout[39]  = hphy_inst_PHYDDIODQDOUT_bus[39];
assign \phy_ddio_dqdout[40]  = hphy_inst_PHYDDIODQDOUT_bus[40];
assign \phy_ddio_dqdout[41]  = hphy_inst_PHYDDIODQDOUT_bus[41];
assign \phy_ddio_dqdout[42]  = hphy_inst_PHYDDIODQDOUT_bus[42];
assign \phy_ddio_dqdout[43]  = hphy_inst_PHYDDIODQDOUT_bus[43];
assign \phy_ddio_dqdout[44]  = hphy_inst_PHYDDIODQDOUT_bus[44];
assign \phy_ddio_dqdout[45]  = hphy_inst_PHYDDIODQDOUT_bus[45];
assign \phy_ddio_dqdout[46]  = hphy_inst_PHYDDIODQDOUT_bus[46];
assign \phy_ddio_dqdout[47]  = hphy_inst_PHYDDIODQDOUT_bus[47];
assign \phy_ddio_dqdout[48]  = hphy_inst_PHYDDIODQDOUT_bus[48];
assign \phy_ddio_dqdout[49]  = hphy_inst_PHYDDIODQDOUT_bus[49];
assign \phy_ddio_dqdout[50]  = hphy_inst_PHYDDIODQDOUT_bus[50];
assign \phy_ddio_dqdout[51]  = hphy_inst_PHYDDIODQDOUT_bus[51];
assign \phy_ddio_dqdout[52]  = hphy_inst_PHYDDIODQDOUT_bus[52];
assign \phy_ddio_dqdout[53]  = hphy_inst_PHYDDIODQDOUT_bus[53];
assign \phy_ddio_dqdout[54]  = hphy_inst_PHYDDIODQDOUT_bus[54];
assign \phy_ddio_dqdout[55]  = hphy_inst_PHYDDIODQDOUT_bus[55];
assign \phy_ddio_dqdout[56]  = hphy_inst_PHYDDIODQDOUT_bus[56];
assign \phy_ddio_dqdout[57]  = hphy_inst_PHYDDIODQDOUT_bus[57];
assign \phy_ddio_dqdout[58]  = hphy_inst_PHYDDIODQDOUT_bus[58];
assign \phy_ddio_dqdout[59]  = hphy_inst_PHYDDIODQDOUT_bus[59];
assign \phy_ddio_dqdout[60]  = hphy_inst_PHYDDIODQDOUT_bus[60];
assign \phy_ddio_dqdout[61]  = hphy_inst_PHYDDIODQDOUT_bus[61];
assign \phy_ddio_dqdout[62]  = hphy_inst_PHYDDIODQDOUT_bus[62];
assign \phy_ddio_dqdout[63]  = hphy_inst_PHYDDIODQDOUT_bus[63];
assign \phy_ddio_dqdout[64]  = hphy_inst_PHYDDIODQDOUT_bus[64];
assign \phy_ddio_dqdout[65]  = hphy_inst_PHYDDIODQDOUT_bus[65];
assign \phy_ddio_dqdout[66]  = hphy_inst_PHYDDIODQDOUT_bus[66];
assign \phy_ddio_dqdout[67]  = hphy_inst_PHYDDIODQDOUT_bus[67];
assign \phy_ddio_dqdout[72]  = hphy_inst_PHYDDIODQDOUT_bus[72];
assign \phy_ddio_dqdout[73]  = hphy_inst_PHYDDIODQDOUT_bus[73];
assign \phy_ddio_dqdout[74]  = hphy_inst_PHYDDIODQDOUT_bus[74];
assign \phy_ddio_dqdout[75]  = hphy_inst_PHYDDIODQDOUT_bus[75];
assign \phy_ddio_dqdout[76]  = hphy_inst_PHYDDIODQDOUT_bus[76];
assign \phy_ddio_dqdout[77]  = hphy_inst_PHYDDIODQDOUT_bus[77];
assign \phy_ddio_dqdout[78]  = hphy_inst_PHYDDIODQDOUT_bus[78];
assign \phy_ddio_dqdout[79]  = hphy_inst_PHYDDIODQDOUT_bus[79];
assign \phy_ddio_dqdout[80]  = hphy_inst_PHYDDIODQDOUT_bus[80];
assign \phy_ddio_dqdout[81]  = hphy_inst_PHYDDIODQDOUT_bus[81];
assign \phy_ddio_dqdout[82]  = hphy_inst_PHYDDIODQDOUT_bus[82];
assign \phy_ddio_dqdout[83]  = hphy_inst_PHYDDIODQDOUT_bus[83];
assign \phy_ddio_dqdout[84]  = hphy_inst_PHYDDIODQDOUT_bus[84];
assign \phy_ddio_dqdout[85]  = hphy_inst_PHYDDIODQDOUT_bus[85];
assign \phy_ddio_dqdout[86]  = hphy_inst_PHYDDIODQDOUT_bus[86];
assign \phy_ddio_dqdout[87]  = hphy_inst_PHYDDIODQDOUT_bus[87];
assign \phy_ddio_dqdout[88]  = hphy_inst_PHYDDIODQDOUT_bus[88];
assign \phy_ddio_dqdout[89]  = hphy_inst_PHYDDIODQDOUT_bus[89];
assign \phy_ddio_dqdout[90]  = hphy_inst_PHYDDIODQDOUT_bus[90];
assign \phy_ddio_dqdout[91]  = hphy_inst_PHYDDIODQDOUT_bus[91];
assign \phy_ddio_dqdout[92]  = hphy_inst_PHYDDIODQDOUT_bus[92];
assign \phy_ddio_dqdout[93]  = hphy_inst_PHYDDIODQDOUT_bus[93];
assign \phy_ddio_dqdout[94]  = hphy_inst_PHYDDIODQDOUT_bus[94];
assign \phy_ddio_dqdout[95]  = hphy_inst_PHYDDIODQDOUT_bus[95];
assign \phy_ddio_dqdout[96]  = hphy_inst_PHYDDIODQDOUT_bus[96];
assign \phy_ddio_dqdout[97]  = hphy_inst_PHYDDIODQDOUT_bus[97];
assign \phy_ddio_dqdout[98]  = hphy_inst_PHYDDIODQDOUT_bus[98];
assign \phy_ddio_dqdout[99]  = hphy_inst_PHYDDIODQDOUT_bus[99];
assign \phy_ddio_dqdout[100]  = hphy_inst_PHYDDIODQDOUT_bus[100];
assign \phy_ddio_dqdout[101]  = hphy_inst_PHYDDIODQDOUT_bus[101];
assign \phy_ddio_dqdout[102]  = hphy_inst_PHYDDIODQDOUT_bus[102];
assign \phy_ddio_dqdout[103]  = hphy_inst_PHYDDIODQDOUT_bus[103];
assign \phy_ddio_dqdout[108]  = hphy_inst_PHYDDIODQDOUT_bus[108];
assign \phy_ddio_dqdout[109]  = hphy_inst_PHYDDIODQDOUT_bus[109];
assign \phy_ddio_dqdout[110]  = hphy_inst_PHYDDIODQDOUT_bus[110];
assign \phy_ddio_dqdout[111]  = hphy_inst_PHYDDIODQDOUT_bus[111];
assign \phy_ddio_dqdout[112]  = hphy_inst_PHYDDIODQDOUT_bus[112];
assign \phy_ddio_dqdout[113]  = hphy_inst_PHYDDIODQDOUT_bus[113];
assign \phy_ddio_dqdout[114]  = hphy_inst_PHYDDIODQDOUT_bus[114];
assign \phy_ddio_dqdout[115]  = hphy_inst_PHYDDIODQDOUT_bus[115];
assign \phy_ddio_dqdout[116]  = hphy_inst_PHYDDIODQDOUT_bus[116];
assign \phy_ddio_dqdout[117]  = hphy_inst_PHYDDIODQDOUT_bus[117];
assign \phy_ddio_dqdout[118]  = hphy_inst_PHYDDIODQDOUT_bus[118];
assign \phy_ddio_dqdout[119]  = hphy_inst_PHYDDIODQDOUT_bus[119];
assign \phy_ddio_dqdout[120]  = hphy_inst_PHYDDIODQDOUT_bus[120];
assign \phy_ddio_dqdout[121]  = hphy_inst_PHYDDIODQDOUT_bus[121];
assign \phy_ddio_dqdout[122]  = hphy_inst_PHYDDIODQDOUT_bus[122];
assign \phy_ddio_dqdout[123]  = hphy_inst_PHYDDIODQDOUT_bus[123];
assign \phy_ddio_dqdout[124]  = hphy_inst_PHYDDIODQDOUT_bus[124];
assign \phy_ddio_dqdout[125]  = hphy_inst_PHYDDIODQDOUT_bus[125];
assign \phy_ddio_dqdout[126]  = hphy_inst_PHYDDIODQDOUT_bus[126];
assign \phy_ddio_dqdout[127]  = hphy_inst_PHYDDIODQDOUT_bus[127];
assign \phy_ddio_dqdout[128]  = hphy_inst_PHYDDIODQDOUT_bus[128];
assign \phy_ddio_dqdout[129]  = hphy_inst_PHYDDIODQDOUT_bus[129];
assign \phy_ddio_dqdout[130]  = hphy_inst_PHYDDIODQDOUT_bus[130];
assign \phy_ddio_dqdout[131]  = hphy_inst_PHYDDIODQDOUT_bus[131];
assign \phy_ddio_dqdout[132]  = hphy_inst_PHYDDIODQDOUT_bus[132];
assign \phy_ddio_dqdout[133]  = hphy_inst_PHYDDIODQDOUT_bus[133];
assign \phy_ddio_dqdout[134]  = hphy_inst_PHYDDIODQDOUT_bus[134];
assign \phy_ddio_dqdout[135]  = hphy_inst_PHYDDIODQDOUT_bus[135];
assign \phy_ddio_dqdout[136]  = hphy_inst_PHYDDIODQDOUT_bus[136];
assign \phy_ddio_dqdout[137]  = hphy_inst_PHYDDIODQDOUT_bus[137];
assign \phy_ddio_dqdout[138]  = hphy_inst_PHYDDIODQDOUT_bus[138];
assign \phy_ddio_dqdout[139]  = hphy_inst_PHYDDIODQDOUT_bus[139];

assign \phy_ddio_dqoe[0]  = hphy_inst_PHYDDIODQOE_bus[0];
assign \phy_ddio_dqoe[1]  = hphy_inst_PHYDDIODQOE_bus[1];
assign \phy_ddio_dqoe[2]  = hphy_inst_PHYDDIODQOE_bus[2];
assign \phy_ddio_dqoe[3]  = hphy_inst_PHYDDIODQOE_bus[3];
assign \phy_ddio_dqoe[4]  = hphy_inst_PHYDDIODQOE_bus[4];
assign \phy_ddio_dqoe[5]  = hphy_inst_PHYDDIODQOE_bus[5];
assign \phy_ddio_dqoe[6]  = hphy_inst_PHYDDIODQOE_bus[6];
assign \phy_ddio_dqoe[7]  = hphy_inst_PHYDDIODQOE_bus[7];
assign \phy_ddio_dqoe[8]  = hphy_inst_PHYDDIODQOE_bus[8];
assign \phy_ddio_dqoe[9]  = hphy_inst_PHYDDIODQOE_bus[9];
assign \phy_ddio_dqoe[10]  = hphy_inst_PHYDDIODQOE_bus[10];
assign \phy_ddio_dqoe[11]  = hphy_inst_PHYDDIODQOE_bus[11];
assign \phy_ddio_dqoe[12]  = hphy_inst_PHYDDIODQOE_bus[12];
assign \phy_ddio_dqoe[13]  = hphy_inst_PHYDDIODQOE_bus[13];
assign \phy_ddio_dqoe[14]  = hphy_inst_PHYDDIODQOE_bus[14];
assign \phy_ddio_dqoe[15]  = hphy_inst_PHYDDIODQOE_bus[15];
assign \phy_ddio_dqoe[18]  = hphy_inst_PHYDDIODQOE_bus[18];
assign \phy_ddio_dqoe[19]  = hphy_inst_PHYDDIODQOE_bus[19];
assign \phy_ddio_dqoe[20]  = hphy_inst_PHYDDIODQOE_bus[20];
assign \phy_ddio_dqoe[21]  = hphy_inst_PHYDDIODQOE_bus[21];
assign \phy_ddio_dqoe[22]  = hphy_inst_PHYDDIODQOE_bus[22];
assign \phy_ddio_dqoe[23]  = hphy_inst_PHYDDIODQOE_bus[23];
assign \phy_ddio_dqoe[24]  = hphy_inst_PHYDDIODQOE_bus[24];
assign \phy_ddio_dqoe[25]  = hphy_inst_PHYDDIODQOE_bus[25];
assign \phy_ddio_dqoe[26]  = hphy_inst_PHYDDIODQOE_bus[26];
assign \phy_ddio_dqoe[27]  = hphy_inst_PHYDDIODQOE_bus[27];
assign \phy_ddio_dqoe[28]  = hphy_inst_PHYDDIODQOE_bus[28];
assign \phy_ddio_dqoe[29]  = hphy_inst_PHYDDIODQOE_bus[29];
assign \phy_ddio_dqoe[30]  = hphy_inst_PHYDDIODQOE_bus[30];
assign \phy_ddio_dqoe[31]  = hphy_inst_PHYDDIODQOE_bus[31];
assign \phy_ddio_dqoe[32]  = hphy_inst_PHYDDIODQOE_bus[32];
assign \phy_ddio_dqoe[33]  = hphy_inst_PHYDDIODQOE_bus[33];
assign \phy_ddio_dqoe[36]  = hphy_inst_PHYDDIODQOE_bus[36];
assign \phy_ddio_dqoe[37]  = hphy_inst_PHYDDIODQOE_bus[37];
assign \phy_ddio_dqoe[38]  = hphy_inst_PHYDDIODQOE_bus[38];
assign \phy_ddio_dqoe[39]  = hphy_inst_PHYDDIODQOE_bus[39];
assign \phy_ddio_dqoe[40]  = hphy_inst_PHYDDIODQOE_bus[40];
assign \phy_ddio_dqoe[41]  = hphy_inst_PHYDDIODQOE_bus[41];
assign \phy_ddio_dqoe[42]  = hphy_inst_PHYDDIODQOE_bus[42];
assign \phy_ddio_dqoe[43]  = hphy_inst_PHYDDIODQOE_bus[43];
assign \phy_ddio_dqoe[44]  = hphy_inst_PHYDDIODQOE_bus[44];
assign \phy_ddio_dqoe[45]  = hphy_inst_PHYDDIODQOE_bus[45];
assign \phy_ddio_dqoe[46]  = hphy_inst_PHYDDIODQOE_bus[46];
assign \phy_ddio_dqoe[47]  = hphy_inst_PHYDDIODQOE_bus[47];
assign \phy_ddio_dqoe[48]  = hphy_inst_PHYDDIODQOE_bus[48];
assign \phy_ddio_dqoe[49]  = hphy_inst_PHYDDIODQOE_bus[49];
assign \phy_ddio_dqoe[50]  = hphy_inst_PHYDDIODQOE_bus[50];
assign \phy_ddio_dqoe[51]  = hphy_inst_PHYDDIODQOE_bus[51];
assign \phy_ddio_dqoe[54]  = hphy_inst_PHYDDIODQOE_bus[54];
assign \phy_ddio_dqoe[55]  = hphy_inst_PHYDDIODQOE_bus[55];
assign \phy_ddio_dqoe[56]  = hphy_inst_PHYDDIODQOE_bus[56];
assign \phy_ddio_dqoe[57]  = hphy_inst_PHYDDIODQOE_bus[57];
assign \phy_ddio_dqoe[58]  = hphy_inst_PHYDDIODQOE_bus[58];
assign \phy_ddio_dqoe[59]  = hphy_inst_PHYDDIODQOE_bus[59];
assign \phy_ddio_dqoe[60]  = hphy_inst_PHYDDIODQOE_bus[60];
assign \phy_ddio_dqoe[61]  = hphy_inst_PHYDDIODQOE_bus[61];
assign \phy_ddio_dqoe[62]  = hphy_inst_PHYDDIODQOE_bus[62];
assign \phy_ddio_dqoe[63]  = hphy_inst_PHYDDIODQOE_bus[63];
assign \phy_ddio_dqoe[64]  = hphy_inst_PHYDDIODQOE_bus[64];
assign \phy_ddio_dqoe[65]  = hphy_inst_PHYDDIODQOE_bus[65];
assign \phy_ddio_dqoe[66]  = hphy_inst_PHYDDIODQOE_bus[66];
assign \phy_ddio_dqoe[67]  = hphy_inst_PHYDDIODQOE_bus[67];
assign \phy_ddio_dqoe[68]  = hphy_inst_PHYDDIODQOE_bus[68];
assign \phy_ddio_dqoe[69]  = hphy_inst_PHYDDIODQOE_bus[69];

assign \phy_ddio_dqs_dout[0]  = hphy_inst_PHYDDIODQSDOUT_bus[0];
assign \phy_ddio_dqs_dout[1]  = hphy_inst_PHYDDIODQSDOUT_bus[1];
assign \phy_ddio_dqs_dout[2]  = hphy_inst_PHYDDIODQSDOUT_bus[2];
assign \phy_ddio_dqs_dout[3]  = hphy_inst_PHYDDIODQSDOUT_bus[3];
assign \phy_ddio_dqs_dout[4]  = hphy_inst_PHYDDIODQSDOUT_bus[4];
assign \phy_ddio_dqs_dout[5]  = hphy_inst_PHYDDIODQSDOUT_bus[5];
assign \phy_ddio_dqs_dout[6]  = hphy_inst_PHYDDIODQSDOUT_bus[6];
assign \phy_ddio_dqs_dout[7]  = hphy_inst_PHYDDIODQSDOUT_bus[7];
assign \phy_ddio_dqs_dout[8]  = hphy_inst_PHYDDIODQSDOUT_bus[8];
assign \phy_ddio_dqs_dout[9]  = hphy_inst_PHYDDIODQSDOUT_bus[9];
assign \phy_ddio_dqs_dout[10]  = hphy_inst_PHYDDIODQSDOUT_bus[10];
assign \phy_ddio_dqs_dout[11]  = hphy_inst_PHYDDIODQSDOUT_bus[11];
assign \phy_ddio_dqs_dout[12]  = hphy_inst_PHYDDIODQSDOUT_bus[12];
assign \phy_ddio_dqs_dout[13]  = hphy_inst_PHYDDIODQSDOUT_bus[13];
assign \phy_ddio_dqs_dout[14]  = hphy_inst_PHYDDIODQSDOUT_bus[14];
assign \phy_ddio_dqs_dout[15]  = hphy_inst_PHYDDIODQSDOUT_bus[15];

assign \phy_ddio_dqslogic_aclr_fifoctrl[0]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[0];
assign \phy_ddio_dqslogic_aclr_fifoctrl[1]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[1];
assign \phy_ddio_dqslogic_aclr_fifoctrl[2]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[2];
assign \phy_ddio_dqslogic_aclr_fifoctrl[3]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[3];

assign \phy_ddio_dqslogic_aclr_pstamble[0]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[0];
assign \phy_ddio_dqslogic_aclr_pstamble[1]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[1];
assign \phy_ddio_dqslogic_aclr_pstamble[2]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[2];
assign \phy_ddio_dqslogic_aclr_pstamble[3]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[3];

assign \phy_ddio_dqslogic_dqsena[0]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[0];
assign \phy_ddio_dqslogic_dqsena[1]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[1];
assign \phy_ddio_dqslogic_dqsena[2]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[2];
assign \phy_ddio_dqslogic_dqsena[3]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[3];
assign \phy_ddio_dqslogic_dqsena[4]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[4];
assign \phy_ddio_dqslogic_dqsena[5]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[5];
assign \phy_ddio_dqslogic_dqsena[6]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[6];
assign \phy_ddio_dqslogic_dqsena[7]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[7];

assign \phy_ddio_dqslogic_fiforeset[0]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[0];
assign \phy_ddio_dqslogic_fiforeset[1]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[1];
assign \phy_ddio_dqslogic_fiforeset[2]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[2];
assign \phy_ddio_dqslogic_fiforeset[3]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[3];

assign \phy_ddio_dqslogic_incrdataen[0]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[0];
assign \phy_ddio_dqslogic_incrdataen[1]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[1];
assign \phy_ddio_dqslogic_incrdataen[2]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[2];
assign \phy_ddio_dqslogic_incrdataen[3]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[3];
assign \phy_ddio_dqslogic_incrdataen[4]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[4];
assign \phy_ddio_dqslogic_incrdataen[5]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[5];
assign \phy_ddio_dqslogic_incrdataen[6]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[6];
assign \phy_ddio_dqslogic_incrdataen[7]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[7];

assign \phy_ddio_dqslogic_incwrptr[0]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[0];
assign \phy_ddio_dqslogic_incwrptr[1]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[1];
assign \phy_ddio_dqslogic_incwrptr[2]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[2];
assign \phy_ddio_dqslogic_incwrptr[3]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[3];
assign \phy_ddio_dqslogic_incwrptr[4]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[4];
assign \phy_ddio_dqslogic_incwrptr[5]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[5];
assign \phy_ddio_dqslogic_incwrptr[6]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[6];
assign \phy_ddio_dqslogic_incwrptr[7]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[7];

assign \phy_ddio_dqslogic_oct[0]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[0];
assign \phy_ddio_dqslogic_oct[1]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[1];
assign \phy_ddio_dqslogic_oct[2]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[2];
assign \phy_ddio_dqslogic_oct[3]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[3];
assign \phy_ddio_dqslogic_oct[4]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[4];
assign \phy_ddio_dqslogic_oct[5]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[5];
assign \phy_ddio_dqslogic_oct[6]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[6];
assign \phy_ddio_dqslogic_oct[7]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[7];

assign \phy_ddio_dqslogic_readlatency[0]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[0];
assign \phy_ddio_dqslogic_readlatency[1]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[1];
assign \phy_ddio_dqslogic_readlatency[2]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[2];
assign \phy_ddio_dqslogic_readlatency[3]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[3];
assign \phy_ddio_dqslogic_readlatency[4]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[4];
assign \phy_ddio_dqslogic_readlatency[5]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[5];
assign \phy_ddio_dqslogic_readlatency[6]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[6];
assign \phy_ddio_dqslogic_readlatency[7]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[7];
assign \phy_ddio_dqslogic_readlatency[8]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[8];
assign \phy_ddio_dqslogic_readlatency[9]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[9];
assign \phy_ddio_dqslogic_readlatency[10]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[10];
assign \phy_ddio_dqslogic_readlatency[11]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[11];
assign \phy_ddio_dqslogic_readlatency[12]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[12];
assign \phy_ddio_dqslogic_readlatency[13]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[13];
assign \phy_ddio_dqslogic_readlatency[14]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[14];
assign \phy_ddio_dqslogic_readlatency[15]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[15];
assign \phy_ddio_dqslogic_readlatency[16]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[16];
assign \phy_ddio_dqslogic_readlatency[17]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[17];
assign \phy_ddio_dqslogic_readlatency[18]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[18];
assign \phy_ddio_dqslogic_readlatency[19]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[19];

assign \phy_ddio_dqs_oe[0]  = hphy_inst_PHYDDIODQSOE_bus[0];
assign \phy_ddio_dqs_oe[1]  = hphy_inst_PHYDDIODQSOE_bus[1];
assign \phy_ddio_dqs_oe[2]  = hphy_inst_PHYDDIODQSOE_bus[2];
assign \phy_ddio_dqs_oe[3]  = hphy_inst_PHYDDIODQSOE_bus[3];
assign \phy_ddio_dqs_oe[4]  = hphy_inst_PHYDDIODQSOE_bus[4];
assign \phy_ddio_dqs_oe[5]  = hphy_inst_PHYDDIODQSOE_bus[5];
assign \phy_ddio_dqs_oe[6]  = hphy_inst_PHYDDIODQSOE_bus[6];
assign \phy_ddio_dqs_oe[7]  = hphy_inst_PHYDDIODQSOE_bus[7];

assign \phy_ddio_odt[0]  = hphy_inst_PHYDDIOODTDOUT_bus[0];
assign \phy_ddio_odt[1]  = hphy_inst_PHYDDIOODTDOUT_bus[1];
assign \phy_ddio_odt[2]  = hphy_inst_PHYDDIOODTDOUT_bus[2];
assign \phy_ddio_odt[3]  = hphy_inst_PHYDDIOODTDOUT_bus[3];

assign \phy_ddio_ras_n[0]  = hphy_inst_PHYDDIORASNDOUT_bus[0];
assign \phy_ddio_ras_n[1]  = hphy_inst_PHYDDIORASNDOUT_bus[1];
assign \phy_ddio_ras_n[2]  = hphy_inst_PHYDDIORASNDOUT_bus[2];
assign \phy_ddio_ras_n[3]  = hphy_inst_PHYDDIORASNDOUT_bus[3];

assign \phy_ddio_reset_n[0]  = hphy_inst_PHYDDIORESETNDOUT_bus[0];
assign \phy_ddio_reset_n[1]  = hphy_inst_PHYDDIORESETNDOUT_bus[1];
assign \phy_ddio_reset_n[2]  = hphy_inst_PHYDDIORESETNDOUT_bus[2];
assign \phy_ddio_reset_n[3]  = hphy_inst_PHYDDIORESETNDOUT_bus[3];

assign \phy_ddio_we_n[0]  = hphy_inst_PHYDDIOWENDOUT_bus[0];
assign \phy_ddio_we_n[1]  = hphy_inst_PHYDDIOWENDOUT_bus[1];
assign \phy_ddio_we_n[2]  = hphy_inst_PHYDDIOWENDOUT_bus[2];
assign \phy_ddio_we_n[3]  = hphy_inst_PHYDDIOWENDOUT_bus[3];

soc_system_hps_sdram_p0_acv_hard_io_pads uio_pads(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(\phy_ddio_address[0] ),
	.phy_ddio_address_1(\phy_ddio_address[1] ),
	.phy_ddio_address_2(\phy_ddio_address[2] ),
	.phy_ddio_address_3(\phy_ddio_address[3] ),
	.phy_ddio_address_4(\phy_ddio_address[4] ),
	.phy_ddio_address_5(\phy_ddio_address[5] ),
	.phy_ddio_address_6(\phy_ddio_address[6] ),
	.phy_ddio_address_7(\phy_ddio_address[7] ),
	.phy_ddio_address_8(\phy_ddio_address[8] ),
	.phy_ddio_address_9(\phy_ddio_address[9] ),
	.phy_ddio_address_10(\phy_ddio_address[10] ),
	.phy_ddio_address_11(\phy_ddio_address[11] ),
	.phy_ddio_address_12(\phy_ddio_address[12] ),
	.phy_ddio_address_13(\phy_ddio_address[13] ),
	.phy_ddio_address_14(\phy_ddio_address[14] ),
	.phy_ddio_address_15(\phy_ddio_address[15] ),
	.phy_ddio_address_16(\phy_ddio_address[16] ),
	.phy_ddio_address_17(\phy_ddio_address[17] ),
	.phy_ddio_address_18(\phy_ddio_address[18] ),
	.phy_ddio_address_19(\phy_ddio_address[19] ),
	.phy_ddio_address_20(\phy_ddio_address[20] ),
	.phy_ddio_address_21(\phy_ddio_address[21] ),
	.phy_ddio_address_22(\phy_ddio_address[22] ),
	.phy_ddio_address_23(\phy_ddio_address[23] ),
	.phy_ddio_address_24(\phy_ddio_address[24] ),
	.phy_ddio_address_25(\phy_ddio_address[25] ),
	.phy_ddio_address_26(\phy_ddio_address[26] ),
	.phy_ddio_address_27(\phy_ddio_address[27] ),
	.phy_ddio_address_28(\phy_ddio_address[28] ),
	.phy_ddio_address_29(\phy_ddio_address[29] ),
	.phy_ddio_address_30(\phy_ddio_address[30] ),
	.phy_ddio_address_31(\phy_ddio_address[31] ),
	.phy_ddio_address_32(\phy_ddio_address[32] ),
	.phy_ddio_address_33(\phy_ddio_address[33] ),
	.phy_ddio_address_34(\phy_ddio_address[34] ),
	.phy_ddio_address_35(\phy_ddio_address[35] ),
	.phy_ddio_address_36(\phy_ddio_address[36] ),
	.phy_ddio_address_37(\phy_ddio_address[37] ),
	.phy_ddio_address_38(\phy_ddio_address[38] ),
	.phy_ddio_address_39(\phy_ddio_address[39] ),
	.phy_ddio_address_40(\phy_ddio_address[40] ),
	.phy_ddio_address_41(\phy_ddio_address[41] ),
	.phy_ddio_address_42(\phy_ddio_address[42] ),
	.phy_ddio_address_43(\phy_ddio_address[43] ),
	.phy_ddio_address_44(\phy_ddio_address[44] ),
	.phy_ddio_address_45(\phy_ddio_address[45] ),
	.phy_ddio_address_46(\phy_ddio_address[46] ),
	.phy_ddio_address_47(\phy_ddio_address[47] ),
	.phy_ddio_address_48(\phy_ddio_address[48] ),
	.phy_ddio_address_49(\phy_ddio_address[49] ),
	.phy_ddio_address_50(\phy_ddio_address[50] ),
	.phy_ddio_address_51(\phy_ddio_address[51] ),
	.phy_ddio_address_52(\phy_ddio_address[52] ),
	.phy_ddio_address_53(\phy_ddio_address[53] ),
	.phy_ddio_address_54(\phy_ddio_address[54] ),
	.phy_ddio_address_55(\phy_ddio_address[55] ),
	.phy_ddio_address_56(\phy_ddio_address[56] ),
	.phy_ddio_address_57(\phy_ddio_address[57] ),
	.phy_ddio_address_58(\phy_ddio_address[58] ),
	.phy_ddio_address_59(\phy_ddio_address[59] ),
	.phy_ddio_bank_0(\phy_ddio_bank[0] ),
	.phy_ddio_bank_1(\phy_ddio_bank[1] ),
	.phy_ddio_bank_2(\phy_ddio_bank[2] ),
	.phy_ddio_bank_3(\phy_ddio_bank[3] ),
	.phy_ddio_bank_4(\phy_ddio_bank[4] ),
	.phy_ddio_bank_5(\phy_ddio_bank[5] ),
	.phy_ddio_bank_6(\phy_ddio_bank[6] ),
	.phy_ddio_bank_7(\phy_ddio_bank[7] ),
	.phy_ddio_bank_8(\phy_ddio_bank[8] ),
	.phy_ddio_bank_9(\phy_ddio_bank[9] ),
	.phy_ddio_bank_10(\phy_ddio_bank[10] ),
	.phy_ddio_bank_11(\phy_ddio_bank[11] ),
	.phy_ddio_cas_n_0(\phy_ddio_cas_n[0] ),
	.phy_ddio_cas_n_1(\phy_ddio_cas_n[1] ),
	.phy_ddio_cas_n_2(\phy_ddio_cas_n[2] ),
	.phy_ddio_cas_n_3(\phy_ddio_cas_n[3] ),
	.phy_ddio_ck_0(\phy_ddio_ck[0] ),
	.phy_ddio_ck_1(\phy_ddio_ck[1] ),
	.phy_ddio_cke_0(\phy_ddio_cke[0] ),
	.phy_ddio_cke_1(\phy_ddio_cke[1] ),
	.phy_ddio_cke_2(\phy_ddio_cke[2] ),
	.phy_ddio_cke_3(\phy_ddio_cke[3] ),
	.phy_ddio_cs_n_0(\phy_ddio_cs_n[0] ),
	.phy_ddio_cs_n_1(\phy_ddio_cs_n[1] ),
	.phy_ddio_cs_n_2(\phy_ddio_cs_n[2] ),
	.phy_ddio_cs_n_3(\phy_ddio_cs_n[3] ),
	.phy_ddio_dmdout_0(\phy_ddio_dmdout[0] ),
	.phy_ddio_dmdout_1(\phy_ddio_dmdout[1] ),
	.phy_ddio_dmdout_2(\phy_ddio_dmdout[2] ),
	.phy_ddio_dmdout_3(\phy_ddio_dmdout[3] ),
	.phy_ddio_dmdout_4(\phy_ddio_dmdout[4] ),
	.phy_ddio_dmdout_5(\phy_ddio_dmdout[5] ),
	.phy_ddio_dmdout_6(\phy_ddio_dmdout[6] ),
	.phy_ddio_dmdout_7(\phy_ddio_dmdout[7] ),
	.phy_ddio_dmdout_8(\phy_ddio_dmdout[8] ),
	.phy_ddio_dmdout_9(\phy_ddio_dmdout[9] ),
	.phy_ddio_dmdout_10(\phy_ddio_dmdout[10] ),
	.phy_ddio_dmdout_11(\phy_ddio_dmdout[11] ),
	.phy_ddio_dmdout_12(\phy_ddio_dmdout[12] ),
	.phy_ddio_dmdout_13(\phy_ddio_dmdout[13] ),
	.phy_ddio_dmdout_14(\phy_ddio_dmdout[14] ),
	.phy_ddio_dmdout_15(\phy_ddio_dmdout[15] ),
	.phy_ddio_dqdout_0(\phy_ddio_dqdout[0] ),
	.phy_ddio_dqdout_1(\phy_ddio_dqdout[1] ),
	.phy_ddio_dqdout_2(\phy_ddio_dqdout[2] ),
	.phy_ddio_dqdout_3(\phy_ddio_dqdout[3] ),
	.phy_ddio_dqdout_4(\phy_ddio_dqdout[4] ),
	.phy_ddio_dqdout_5(\phy_ddio_dqdout[5] ),
	.phy_ddio_dqdout_6(\phy_ddio_dqdout[6] ),
	.phy_ddio_dqdout_7(\phy_ddio_dqdout[7] ),
	.phy_ddio_dqdout_8(\phy_ddio_dqdout[8] ),
	.phy_ddio_dqdout_9(\phy_ddio_dqdout[9] ),
	.phy_ddio_dqdout_10(\phy_ddio_dqdout[10] ),
	.phy_ddio_dqdout_11(\phy_ddio_dqdout[11] ),
	.phy_ddio_dqdout_12(\phy_ddio_dqdout[12] ),
	.phy_ddio_dqdout_13(\phy_ddio_dqdout[13] ),
	.phy_ddio_dqdout_14(\phy_ddio_dqdout[14] ),
	.phy_ddio_dqdout_15(\phy_ddio_dqdout[15] ),
	.phy_ddio_dqdout_16(\phy_ddio_dqdout[16] ),
	.phy_ddio_dqdout_17(\phy_ddio_dqdout[17] ),
	.phy_ddio_dqdout_18(\phy_ddio_dqdout[18] ),
	.phy_ddio_dqdout_19(\phy_ddio_dqdout[19] ),
	.phy_ddio_dqdout_20(\phy_ddio_dqdout[20] ),
	.phy_ddio_dqdout_21(\phy_ddio_dqdout[21] ),
	.phy_ddio_dqdout_22(\phy_ddio_dqdout[22] ),
	.phy_ddio_dqdout_23(\phy_ddio_dqdout[23] ),
	.phy_ddio_dqdout_24(\phy_ddio_dqdout[24] ),
	.phy_ddio_dqdout_25(\phy_ddio_dqdout[25] ),
	.phy_ddio_dqdout_26(\phy_ddio_dqdout[26] ),
	.phy_ddio_dqdout_27(\phy_ddio_dqdout[27] ),
	.phy_ddio_dqdout_28(\phy_ddio_dqdout[28] ),
	.phy_ddio_dqdout_29(\phy_ddio_dqdout[29] ),
	.phy_ddio_dqdout_30(\phy_ddio_dqdout[30] ),
	.phy_ddio_dqdout_31(\phy_ddio_dqdout[31] ),
	.phy_ddio_dqdout_36(\phy_ddio_dqdout[36] ),
	.phy_ddio_dqdout_37(\phy_ddio_dqdout[37] ),
	.phy_ddio_dqdout_38(\phy_ddio_dqdout[38] ),
	.phy_ddio_dqdout_39(\phy_ddio_dqdout[39] ),
	.phy_ddio_dqdout_40(\phy_ddio_dqdout[40] ),
	.phy_ddio_dqdout_41(\phy_ddio_dqdout[41] ),
	.phy_ddio_dqdout_42(\phy_ddio_dqdout[42] ),
	.phy_ddio_dqdout_43(\phy_ddio_dqdout[43] ),
	.phy_ddio_dqdout_44(\phy_ddio_dqdout[44] ),
	.phy_ddio_dqdout_45(\phy_ddio_dqdout[45] ),
	.phy_ddio_dqdout_46(\phy_ddio_dqdout[46] ),
	.phy_ddio_dqdout_47(\phy_ddio_dqdout[47] ),
	.phy_ddio_dqdout_48(\phy_ddio_dqdout[48] ),
	.phy_ddio_dqdout_49(\phy_ddio_dqdout[49] ),
	.phy_ddio_dqdout_50(\phy_ddio_dqdout[50] ),
	.phy_ddio_dqdout_51(\phy_ddio_dqdout[51] ),
	.phy_ddio_dqdout_52(\phy_ddio_dqdout[52] ),
	.phy_ddio_dqdout_53(\phy_ddio_dqdout[53] ),
	.phy_ddio_dqdout_54(\phy_ddio_dqdout[54] ),
	.phy_ddio_dqdout_55(\phy_ddio_dqdout[55] ),
	.phy_ddio_dqdout_56(\phy_ddio_dqdout[56] ),
	.phy_ddio_dqdout_57(\phy_ddio_dqdout[57] ),
	.phy_ddio_dqdout_58(\phy_ddio_dqdout[58] ),
	.phy_ddio_dqdout_59(\phy_ddio_dqdout[59] ),
	.phy_ddio_dqdout_60(\phy_ddio_dqdout[60] ),
	.phy_ddio_dqdout_61(\phy_ddio_dqdout[61] ),
	.phy_ddio_dqdout_62(\phy_ddio_dqdout[62] ),
	.phy_ddio_dqdout_63(\phy_ddio_dqdout[63] ),
	.phy_ddio_dqdout_64(\phy_ddio_dqdout[64] ),
	.phy_ddio_dqdout_65(\phy_ddio_dqdout[65] ),
	.phy_ddio_dqdout_66(\phy_ddio_dqdout[66] ),
	.phy_ddio_dqdout_67(\phy_ddio_dqdout[67] ),
	.phy_ddio_dqdout_72(\phy_ddio_dqdout[72] ),
	.phy_ddio_dqdout_73(\phy_ddio_dqdout[73] ),
	.phy_ddio_dqdout_74(\phy_ddio_dqdout[74] ),
	.phy_ddio_dqdout_75(\phy_ddio_dqdout[75] ),
	.phy_ddio_dqdout_76(\phy_ddio_dqdout[76] ),
	.phy_ddio_dqdout_77(\phy_ddio_dqdout[77] ),
	.phy_ddio_dqdout_78(\phy_ddio_dqdout[78] ),
	.phy_ddio_dqdout_79(\phy_ddio_dqdout[79] ),
	.phy_ddio_dqdout_80(\phy_ddio_dqdout[80] ),
	.phy_ddio_dqdout_81(\phy_ddio_dqdout[81] ),
	.phy_ddio_dqdout_82(\phy_ddio_dqdout[82] ),
	.phy_ddio_dqdout_83(\phy_ddio_dqdout[83] ),
	.phy_ddio_dqdout_84(\phy_ddio_dqdout[84] ),
	.phy_ddio_dqdout_85(\phy_ddio_dqdout[85] ),
	.phy_ddio_dqdout_86(\phy_ddio_dqdout[86] ),
	.phy_ddio_dqdout_87(\phy_ddio_dqdout[87] ),
	.phy_ddio_dqdout_88(\phy_ddio_dqdout[88] ),
	.phy_ddio_dqdout_89(\phy_ddio_dqdout[89] ),
	.phy_ddio_dqdout_90(\phy_ddio_dqdout[90] ),
	.phy_ddio_dqdout_91(\phy_ddio_dqdout[91] ),
	.phy_ddio_dqdout_92(\phy_ddio_dqdout[92] ),
	.phy_ddio_dqdout_93(\phy_ddio_dqdout[93] ),
	.phy_ddio_dqdout_94(\phy_ddio_dqdout[94] ),
	.phy_ddio_dqdout_95(\phy_ddio_dqdout[95] ),
	.phy_ddio_dqdout_96(\phy_ddio_dqdout[96] ),
	.phy_ddio_dqdout_97(\phy_ddio_dqdout[97] ),
	.phy_ddio_dqdout_98(\phy_ddio_dqdout[98] ),
	.phy_ddio_dqdout_99(\phy_ddio_dqdout[99] ),
	.phy_ddio_dqdout_100(\phy_ddio_dqdout[100] ),
	.phy_ddio_dqdout_101(\phy_ddio_dqdout[101] ),
	.phy_ddio_dqdout_102(\phy_ddio_dqdout[102] ),
	.phy_ddio_dqdout_103(\phy_ddio_dqdout[103] ),
	.phy_ddio_dqdout_108(\phy_ddio_dqdout[108] ),
	.phy_ddio_dqdout_109(\phy_ddio_dqdout[109] ),
	.phy_ddio_dqdout_110(\phy_ddio_dqdout[110] ),
	.phy_ddio_dqdout_111(\phy_ddio_dqdout[111] ),
	.phy_ddio_dqdout_112(\phy_ddio_dqdout[112] ),
	.phy_ddio_dqdout_113(\phy_ddio_dqdout[113] ),
	.phy_ddio_dqdout_114(\phy_ddio_dqdout[114] ),
	.phy_ddio_dqdout_115(\phy_ddio_dqdout[115] ),
	.phy_ddio_dqdout_116(\phy_ddio_dqdout[116] ),
	.phy_ddio_dqdout_117(\phy_ddio_dqdout[117] ),
	.phy_ddio_dqdout_118(\phy_ddio_dqdout[118] ),
	.phy_ddio_dqdout_119(\phy_ddio_dqdout[119] ),
	.phy_ddio_dqdout_120(\phy_ddio_dqdout[120] ),
	.phy_ddio_dqdout_121(\phy_ddio_dqdout[121] ),
	.phy_ddio_dqdout_122(\phy_ddio_dqdout[122] ),
	.phy_ddio_dqdout_123(\phy_ddio_dqdout[123] ),
	.phy_ddio_dqdout_124(\phy_ddio_dqdout[124] ),
	.phy_ddio_dqdout_125(\phy_ddio_dqdout[125] ),
	.phy_ddio_dqdout_126(\phy_ddio_dqdout[126] ),
	.phy_ddio_dqdout_127(\phy_ddio_dqdout[127] ),
	.phy_ddio_dqdout_128(\phy_ddio_dqdout[128] ),
	.phy_ddio_dqdout_129(\phy_ddio_dqdout[129] ),
	.phy_ddio_dqdout_130(\phy_ddio_dqdout[130] ),
	.phy_ddio_dqdout_131(\phy_ddio_dqdout[131] ),
	.phy_ddio_dqdout_132(\phy_ddio_dqdout[132] ),
	.phy_ddio_dqdout_133(\phy_ddio_dqdout[133] ),
	.phy_ddio_dqdout_134(\phy_ddio_dqdout[134] ),
	.phy_ddio_dqdout_135(\phy_ddio_dqdout[135] ),
	.phy_ddio_dqdout_136(\phy_ddio_dqdout[136] ),
	.phy_ddio_dqdout_137(\phy_ddio_dqdout[137] ),
	.phy_ddio_dqdout_138(\phy_ddio_dqdout[138] ),
	.phy_ddio_dqdout_139(\phy_ddio_dqdout[139] ),
	.phy_ddio_dqoe_0(\phy_ddio_dqoe[0] ),
	.phy_ddio_dqoe_1(\phy_ddio_dqoe[1] ),
	.phy_ddio_dqoe_2(\phy_ddio_dqoe[2] ),
	.phy_ddio_dqoe_3(\phy_ddio_dqoe[3] ),
	.phy_ddio_dqoe_4(\phy_ddio_dqoe[4] ),
	.phy_ddio_dqoe_5(\phy_ddio_dqoe[5] ),
	.phy_ddio_dqoe_6(\phy_ddio_dqoe[6] ),
	.phy_ddio_dqoe_7(\phy_ddio_dqoe[7] ),
	.phy_ddio_dqoe_8(\phy_ddio_dqoe[8] ),
	.phy_ddio_dqoe_9(\phy_ddio_dqoe[9] ),
	.phy_ddio_dqoe_10(\phy_ddio_dqoe[10] ),
	.phy_ddio_dqoe_11(\phy_ddio_dqoe[11] ),
	.phy_ddio_dqoe_12(\phy_ddio_dqoe[12] ),
	.phy_ddio_dqoe_13(\phy_ddio_dqoe[13] ),
	.phy_ddio_dqoe_14(\phy_ddio_dqoe[14] ),
	.phy_ddio_dqoe_15(\phy_ddio_dqoe[15] ),
	.phy_ddio_dqoe_18(\phy_ddio_dqoe[18] ),
	.phy_ddio_dqoe_19(\phy_ddio_dqoe[19] ),
	.phy_ddio_dqoe_20(\phy_ddio_dqoe[20] ),
	.phy_ddio_dqoe_21(\phy_ddio_dqoe[21] ),
	.phy_ddio_dqoe_22(\phy_ddio_dqoe[22] ),
	.phy_ddio_dqoe_23(\phy_ddio_dqoe[23] ),
	.phy_ddio_dqoe_24(\phy_ddio_dqoe[24] ),
	.phy_ddio_dqoe_25(\phy_ddio_dqoe[25] ),
	.phy_ddio_dqoe_26(\phy_ddio_dqoe[26] ),
	.phy_ddio_dqoe_27(\phy_ddio_dqoe[27] ),
	.phy_ddio_dqoe_28(\phy_ddio_dqoe[28] ),
	.phy_ddio_dqoe_29(\phy_ddio_dqoe[29] ),
	.phy_ddio_dqoe_30(\phy_ddio_dqoe[30] ),
	.phy_ddio_dqoe_31(\phy_ddio_dqoe[31] ),
	.phy_ddio_dqoe_32(\phy_ddio_dqoe[32] ),
	.phy_ddio_dqoe_33(\phy_ddio_dqoe[33] ),
	.phy_ddio_dqoe_36(\phy_ddio_dqoe[36] ),
	.phy_ddio_dqoe_37(\phy_ddio_dqoe[37] ),
	.phy_ddio_dqoe_38(\phy_ddio_dqoe[38] ),
	.phy_ddio_dqoe_39(\phy_ddio_dqoe[39] ),
	.phy_ddio_dqoe_40(\phy_ddio_dqoe[40] ),
	.phy_ddio_dqoe_41(\phy_ddio_dqoe[41] ),
	.phy_ddio_dqoe_42(\phy_ddio_dqoe[42] ),
	.phy_ddio_dqoe_43(\phy_ddio_dqoe[43] ),
	.phy_ddio_dqoe_44(\phy_ddio_dqoe[44] ),
	.phy_ddio_dqoe_45(\phy_ddio_dqoe[45] ),
	.phy_ddio_dqoe_46(\phy_ddio_dqoe[46] ),
	.phy_ddio_dqoe_47(\phy_ddio_dqoe[47] ),
	.phy_ddio_dqoe_48(\phy_ddio_dqoe[48] ),
	.phy_ddio_dqoe_49(\phy_ddio_dqoe[49] ),
	.phy_ddio_dqoe_50(\phy_ddio_dqoe[50] ),
	.phy_ddio_dqoe_51(\phy_ddio_dqoe[51] ),
	.phy_ddio_dqoe_54(\phy_ddio_dqoe[54] ),
	.phy_ddio_dqoe_55(\phy_ddio_dqoe[55] ),
	.phy_ddio_dqoe_56(\phy_ddio_dqoe[56] ),
	.phy_ddio_dqoe_57(\phy_ddio_dqoe[57] ),
	.phy_ddio_dqoe_58(\phy_ddio_dqoe[58] ),
	.phy_ddio_dqoe_59(\phy_ddio_dqoe[59] ),
	.phy_ddio_dqoe_60(\phy_ddio_dqoe[60] ),
	.phy_ddio_dqoe_61(\phy_ddio_dqoe[61] ),
	.phy_ddio_dqoe_62(\phy_ddio_dqoe[62] ),
	.phy_ddio_dqoe_63(\phy_ddio_dqoe[63] ),
	.phy_ddio_dqoe_64(\phy_ddio_dqoe[64] ),
	.phy_ddio_dqoe_65(\phy_ddio_dqoe[65] ),
	.phy_ddio_dqoe_66(\phy_ddio_dqoe[66] ),
	.phy_ddio_dqoe_67(\phy_ddio_dqoe[67] ),
	.phy_ddio_dqoe_68(\phy_ddio_dqoe[68] ),
	.phy_ddio_dqoe_69(\phy_ddio_dqoe[69] ),
	.phy_ddio_dqs_dout_0(\phy_ddio_dqs_dout[0] ),
	.phy_ddio_dqs_dout_1(\phy_ddio_dqs_dout[1] ),
	.phy_ddio_dqs_dout_2(\phy_ddio_dqs_dout[2] ),
	.phy_ddio_dqs_dout_3(\phy_ddio_dqs_dout[3] ),
	.phy_ddio_dqs_dout_4(\phy_ddio_dqs_dout[4] ),
	.phy_ddio_dqs_dout_5(\phy_ddio_dqs_dout[5] ),
	.phy_ddio_dqs_dout_6(\phy_ddio_dqs_dout[6] ),
	.phy_ddio_dqs_dout_7(\phy_ddio_dqs_dout[7] ),
	.phy_ddio_dqs_dout_8(\phy_ddio_dqs_dout[8] ),
	.phy_ddio_dqs_dout_9(\phy_ddio_dqs_dout[9] ),
	.phy_ddio_dqs_dout_10(\phy_ddio_dqs_dout[10] ),
	.phy_ddio_dqs_dout_11(\phy_ddio_dqs_dout[11] ),
	.phy_ddio_dqs_dout_12(\phy_ddio_dqs_dout[12] ),
	.phy_ddio_dqs_dout_13(\phy_ddio_dqs_dout[13] ),
	.phy_ddio_dqs_dout_14(\phy_ddio_dqs_dout[14] ),
	.phy_ddio_dqs_dout_15(\phy_ddio_dqs_dout[15] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(\phy_ddio_dqslogic_aclr_fifoctrl[0] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(\phy_ddio_dqslogic_aclr_fifoctrl[1] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(\phy_ddio_dqslogic_aclr_fifoctrl[2] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(\phy_ddio_dqslogic_aclr_fifoctrl[3] ),
	.phy_ddio_dqslogic_aclr_pstamble_0(\phy_ddio_dqslogic_aclr_pstamble[0] ),
	.phy_ddio_dqslogic_aclr_pstamble_1(\phy_ddio_dqslogic_aclr_pstamble[1] ),
	.phy_ddio_dqslogic_aclr_pstamble_2(\phy_ddio_dqslogic_aclr_pstamble[2] ),
	.phy_ddio_dqslogic_aclr_pstamble_3(\phy_ddio_dqslogic_aclr_pstamble[3] ),
	.phy_ddio_dqslogic_dqsena_0(\phy_ddio_dqslogic_dqsena[0] ),
	.phy_ddio_dqslogic_dqsena_1(\phy_ddio_dqslogic_dqsena[1] ),
	.phy_ddio_dqslogic_dqsena_2(\phy_ddio_dqslogic_dqsena[2] ),
	.phy_ddio_dqslogic_dqsena_3(\phy_ddio_dqslogic_dqsena[3] ),
	.phy_ddio_dqslogic_dqsena_4(\phy_ddio_dqslogic_dqsena[4] ),
	.phy_ddio_dqslogic_dqsena_5(\phy_ddio_dqslogic_dqsena[5] ),
	.phy_ddio_dqslogic_dqsena_6(\phy_ddio_dqslogic_dqsena[6] ),
	.phy_ddio_dqslogic_dqsena_7(\phy_ddio_dqslogic_dqsena[7] ),
	.phy_ddio_dqslogic_fiforeset_0(\phy_ddio_dqslogic_fiforeset[0] ),
	.phy_ddio_dqslogic_fiforeset_1(\phy_ddio_dqslogic_fiforeset[1] ),
	.phy_ddio_dqslogic_fiforeset_2(\phy_ddio_dqslogic_fiforeset[2] ),
	.phy_ddio_dqslogic_fiforeset_3(\phy_ddio_dqslogic_fiforeset[3] ),
	.phy_ddio_dqslogic_incrdataen_0(\phy_ddio_dqslogic_incrdataen[0] ),
	.phy_ddio_dqslogic_incrdataen_1(\phy_ddio_dqslogic_incrdataen[1] ),
	.phy_ddio_dqslogic_incrdataen_2(\phy_ddio_dqslogic_incrdataen[2] ),
	.phy_ddio_dqslogic_incrdataen_3(\phy_ddio_dqslogic_incrdataen[3] ),
	.phy_ddio_dqslogic_incrdataen_4(\phy_ddio_dqslogic_incrdataen[4] ),
	.phy_ddio_dqslogic_incrdataen_5(\phy_ddio_dqslogic_incrdataen[5] ),
	.phy_ddio_dqslogic_incrdataen_6(\phy_ddio_dqslogic_incrdataen[6] ),
	.phy_ddio_dqslogic_incrdataen_7(\phy_ddio_dqslogic_incrdataen[7] ),
	.phy_ddio_dqslogic_incwrptr_0(\phy_ddio_dqslogic_incwrptr[0] ),
	.phy_ddio_dqslogic_incwrptr_1(\phy_ddio_dqslogic_incwrptr[1] ),
	.phy_ddio_dqslogic_incwrptr_2(\phy_ddio_dqslogic_incwrptr[2] ),
	.phy_ddio_dqslogic_incwrptr_3(\phy_ddio_dqslogic_incwrptr[3] ),
	.phy_ddio_dqslogic_incwrptr_4(\phy_ddio_dqslogic_incwrptr[4] ),
	.phy_ddio_dqslogic_incwrptr_5(\phy_ddio_dqslogic_incwrptr[5] ),
	.phy_ddio_dqslogic_incwrptr_6(\phy_ddio_dqslogic_incwrptr[6] ),
	.phy_ddio_dqslogic_incwrptr_7(\phy_ddio_dqslogic_incwrptr[7] ),
	.phy_ddio_dqslogic_oct_0(\phy_ddio_dqslogic_oct[0] ),
	.phy_ddio_dqslogic_oct_1(\phy_ddio_dqslogic_oct[1] ),
	.phy_ddio_dqslogic_oct_2(\phy_ddio_dqslogic_oct[2] ),
	.phy_ddio_dqslogic_oct_3(\phy_ddio_dqslogic_oct[3] ),
	.phy_ddio_dqslogic_oct_4(\phy_ddio_dqslogic_oct[4] ),
	.phy_ddio_dqslogic_oct_5(\phy_ddio_dqslogic_oct[5] ),
	.phy_ddio_dqslogic_oct_6(\phy_ddio_dqslogic_oct[6] ),
	.phy_ddio_dqslogic_oct_7(\phy_ddio_dqslogic_oct[7] ),
	.phy_ddio_dqslogic_readlatency_0(\phy_ddio_dqslogic_readlatency[0] ),
	.phy_ddio_dqslogic_readlatency_1(\phy_ddio_dqslogic_readlatency[1] ),
	.phy_ddio_dqslogic_readlatency_2(\phy_ddio_dqslogic_readlatency[2] ),
	.phy_ddio_dqslogic_readlatency_3(\phy_ddio_dqslogic_readlatency[3] ),
	.phy_ddio_dqslogic_readlatency_4(\phy_ddio_dqslogic_readlatency[4] ),
	.phy_ddio_dqslogic_readlatency_5(\phy_ddio_dqslogic_readlatency[5] ),
	.phy_ddio_dqslogic_readlatency_6(\phy_ddio_dqslogic_readlatency[6] ),
	.phy_ddio_dqslogic_readlatency_7(\phy_ddio_dqslogic_readlatency[7] ),
	.phy_ddio_dqslogic_readlatency_8(\phy_ddio_dqslogic_readlatency[8] ),
	.phy_ddio_dqslogic_readlatency_9(\phy_ddio_dqslogic_readlatency[9] ),
	.phy_ddio_dqslogic_readlatency_10(\phy_ddio_dqslogic_readlatency[10] ),
	.phy_ddio_dqslogic_readlatency_11(\phy_ddio_dqslogic_readlatency[11] ),
	.phy_ddio_dqslogic_readlatency_12(\phy_ddio_dqslogic_readlatency[12] ),
	.phy_ddio_dqslogic_readlatency_13(\phy_ddio_dqslogic_readlatency[13] ),
	.phy_ddio_dqslogic_readlatency_14(\phy_ddio_dqslogic_readlatency[14] ),
	.phy_ddio_dqslogic_readlatency_15(\phy_ddio_dqslogic_readlatency[15] ),
	.phy_ddio_dqslogic_readlatency_16(\phy_ddio_dqslogic_readlatency[16] ),
	.phy_ddio_dqslogic_readlatency_17(\phy_ddio_dqslogic_readlatency[17] ),
	.phy_ddio_dqslogic_readlatency_18(\phy_ddio_dqslogic_readlatency[18] ),
	.phy_ddio_dqslogic_readlatency_19(\phy_ddio_dqslogic_readlatency[19] ),
	.phy_ddio_dqs_oe_0(\phy_ddio_dqs_oe[0] ),
	.phy_ddio_dqs_oe_1(\phy_ddio_dqs_oe[1] ),
	.phy_ddio_dqs_oe_2(\phy_ddio_dqs_oe[2] ),
	.phy_ddio_dqs_oe_3(\phy_ddio_dqs_oe[3] ),
	.phy_ddio_dqs_oe_4(\phy_ddio_dqs_oe[4] ),
	.phy_ddio_dqs_oe_5(\phy_ddio_dqs_oe[5] ),
	.phy_ddio_dqs_oe_6(\phy_ddio_dqs_oe[6] ),
	.phy_ddio_dqs_oe_7(\phy_ddio_dqs_oe[7] ),
	.phy_ddio_odt_0(\phy_ddio_odt[0] ),
	.phy_ddio_odt_1(\phy_ddio_odt[1] ),
	.phy_ddio_odt_2(\phy_ddio_odt[2] ),
	.phy_ddio_odt_3(\phy_ddio_odt[3] ),
	.phy_ddio_ras_n_0(\phy_ddio_ras_n[0] ),
	.phy_ddio_ras_n_1(\phy_ddio_ras_n[1] ),
	.phy_ddio_ras_n_2(\phy_ddio_ras_n[2] ),
	.phy_ddio_ras_n_3(\phy_ddio_ras_n[3] ),
	.phy_ddio_reset_n_0(\phy_ddio_reset_n[0] ),
	.phy_ddio_reset_n_1(\phy_ddio_reset_n[1] ),
	.phy_ddio_reset_n_2(\phy_ddio_reset_n[2] ),
	.phy_ddio_reset_n_3(\phy_ddio_reset_n[3] ),
	.phy_ddio_we_n_0(\phy_ddio_we_n[0] ),
	.phy_ddio_we_n_1(\phy_ddio_we_n[1] ),
	.phy_ddio_we_n_2(\phy_ddio_we_n[2] ),
	.phy_ddio_we_n_3(\phy_ddio_we_n[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.ddio_phy_dqslogic_rdatavalid({ddio_phy_dqslogic_rdatavalid_unconnected_wire_4,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

soc_system_hps_sdram_p0_acv_ldc_25 memphy_ldc(
	.pll_hr_clk(afi_clk),
	.pll_dqs_clk(afi_clk),
	.adc_clk(leveled_dqs_clocks_0),
	.avl_clk(\memphy_ldc|leveled_hr_clocks[0] ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_mem_phy hphy_inst(
	.aficasn(afi_cas_n[0]),
	.afimemclkdisable(afi_mem_clk_disable[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.avlread(gnd),
	.avlresetn(gnd),
	.avlwrite(gnd),
	.globalresetn(gnd),
	.iointcasnaclr(gnd),
	.iointrasnaclr(gnd),
	.iointresetnaclr(gnd),
	.iointwenaclr(gnd),
	.plladdrcmdclk(!leveled_dqs_clocks_0),
	.pllaficlk(leveled_dqs_clocks_0),
	.pllavlclk(\memphy_ldc|leveled_hr_clocks[0] ),
	.plllocked(gnd),
	.scanen(gnd),
	.softresetn(gnd),
	.afiaddr({afi_addr[19],afi_addr[18],afi_addr[17],afi_addr[16],afi_addr[15],afi_addr[14],afi_addr[13],afi_addr[12],afi_addr[11],afi_addr[10],afi_addr[9],afi_addr[8],afi_addr[7],afi_addr[6],afi_addr[5],afi_addr[4],afi_addr[3],afi_addr[2],afi_addr[1],afi_addr[0]}),
	.afiba({afi_ba[2],afi_ba[1],afi_ba[0]}),
	.aficke({afi_cke[1],afi_cke[0]}),
	.aficsn({afi_cs_n[1],afi_cs_n[0]}),
	.afidm({afi_dm[9],afi_dm[8],afi_dm[7],afi_dm[6],afi_dm[5],afi_dm[4],afi_dm[3],afi_dm[2],afi_dm[1],afi_dm[0]}),
	.afidqsburst({afi_dqs_burst[4],afi_dqs_burst[3],afi_dqs_burst[2],afi_dqs_burst[1],afi_dqs_burst[0]}),
	.afiodt({afi_odt[1],afi_odt[0]}),
	.afirdataen({afi_rdata_en[4],afi_rdata_en[3],afi_rdata_en[2],afi_rdata_en[1],afi_rdata_en[0]}),
	.afirdataenfull({afi_rdata_en_full[4],afi_rdata_en_full[3],afi_rdata_en_full[2],afi_rdata_en_full[1],afi_rdata_en_full[0]}),
	.afiwdata({afi_wdata[79],afi_wdata[78],afi_wdata[77],afi_wdata[76],afi_wdata[75],afi_wdata[74],afi_wdata[73],afi_wdata[72],afi_wdata[71],afi_wdata[70],afi_wdata[69],afi_wdata[68],afi_wdata[67],afi_wdata[66],afi_wdata[65],afi_wdata[64],afi_wdata[63],afi_wdata[62],afi_wdata[61],afi_wdata[60],afi_wdata[59],afi_wdata[58],afi_wdata[57],afi_wdata[56],afi_wdata[55],afi_wdata[54],afi_wdata[53],afi_wdata[52],
afi_wdata[51],afi_wdata[50],afi_wdata[49],afi_wdata[48],afi_wdata[47],afi_wdata[46],afi_wdata[45],afi_wdata[44],afi_wdata[43],afi_wdata[42],afi_wdata[41],afi_wdata[40],afi_wdata[39],afi_wdata[38],afi_wdata[37],afi_wdata[36],afi_wdata[35],afi_wdata[34],afi_wdata[33],afi_wdata[32],afi_wdata[31],afi_wdata[30],afi_wdata[29],afi_wdata[28],afi_wdata[27],afi_wdata[26],afi_wdata[25],afi_wdata[24],
afi_wdata[23],afi_wdata[22],afi_wdata[21],afi_wdata[20],afi_wdata[19],afi_wdata[18],afi_wdata[17],afi_wdata[16],afi_wdata[15],afi_wdata[14],afi_wdata[13],afi_wdata[12],afi_wdata[11],afi_wdata[10],afi_wdata[9],afi_wdata[8],afi_wdata[7],afi_wdata[6],afi_wdata[5],afi_wdata[4],afi_wdata[3],afi_wdata[2],afi_wdata[1],afi_wdata[0]}),
	.afiwdatavalid({afi_wdata_valid[4],afi_wdata_valid[3],afi_wdata_valid[2],afi_wdata_valid[1],afi_wdata_valid[0]}),
	.avladdress({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.avlwritedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfgaddlat({gnd,gnd,gnd,cfg_addlat[4],cfg_addlat[3],cfg_addlat[2],cfg_addlat[1],cfg_addlat[0]}),
	.cfgbankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth[2],cfg_bankaddrwidth[1],cfg_bankaddrwidth[0]}),
	.cfgcaswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat[3],cfg_caswrlat[2],cfg_caswrlat[1],cfg_caswrlat[0]}),
	.cfgcoladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth[4],cfg_coladdrwidth[3],cfg_coladdrwidth[2],cfg_coladdrwidth[1],cfg_coladdrwidth[0]}),
	.cfgcsaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth[2],cfg_csaddrwidth[1],cfg_csaddrwidth[0]}),
	.cfgdevicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth[3],cfg_devicewidth[2],cfg_devicewidth[1],cfg_devicewidth[0]}),
	.cfgdramconfig({gnd,gnd,gnd,cfg_dramconfig[20],cfg_dramconfig[19],cfg_dramconfig[18],cfg_dramconfig[17],cfg_dramconfig[16],cfg_dramconfig[15],cfg_dramconfig[14],cfg_dramconfig[13],cfg_dramconfig[12],cfg_dramconfig[11],cfg_dramconfig[10],cfg_dramconfig[9],cfg_dramconfig[8],cfg_dramconfig[7],cfg_dramconfig[6],cfg_dramconfig[5],cfg_dramconfig[4],
cfg_dramconfig[3],cfg_dramconfig[2],cfg_dramconfig[1],cfg_dramconfig[0]}),
	.cfginterfacewidth({cfg_interfacewidth[7],cfg_interfacewidth[6],cfg_interfacewidth[5],cfg_interfacewidth[4],cfg_interfacewidth[3],cfg_interfacewidth[2],cfg_interfacewidth[1],cfg_interfacewidth[0]}),
	.cfgrowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth[4],cfg_rowaddrwidth[3],cfg_rowaddrwidth[2],cfg_rowaddrwidth[1],cfg_rowaddrwidth[0]}),
	.cfgtcl({gnd,gnd,gnd,cfg_tcl[4],cfg_tcl[3],cfg_tcl[2],cfg_tcl[1],cfg_tcl[0]}),
	.cfgtmrd({gnd,gnd,gnd,gnd,cfg_tmrd[3],cfg_tmrd[2],cfg_tmrd[1],cfg_tmrd[0]}),
	.cfgtrefi({gnd,gnd,gnd,cfg_trefi[12],cfg_trefi[11],cfg_trefi[10],cfg_trefi[9],cfg_trefi[8],cfg_trefi[7],cfg_trefi[6],cfg_trefi[5],cfg_trefi[4],cfg_trefi[3],cfg_trefi[2],cfg_trefi[1],cfg_trefi[0]}),
	.cfgtrfc({cfg_trfc[7],cfg_trfc[6],cfg_trfc[5],cfg_trfc[4],cfg_trfc[3],cfg_trfc[2],cfg_trfc[1],cfg_trfc[0]}),
	.cfgtwr({gnd,gnd,gnd,gnd,cfg_twr[3],cfg_twr[2],cfg_twr[1],cfg_twr[0]}),
	.ddiophydqdin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] }),
	.ddiophydqslogicrdatavalid({vcc,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.iointaddraclr(16'b0000000000000000),
	.iointaddrdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointbaaclr(3'b000),
	.iointbadout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointcasndout({gnd,gnd,gnd,gnd}),
	.iointckdout({gnd,gnd,gnd,gnd}),
	.iointckeaclr(2'b00),
	.iointckedout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointckndout({gnd,gnd,gnd,gnd}),
	.iointcsnaclr(2'b00),
	.iointcsndout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdmdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iointdqsbdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsboe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicaclrfifoctrl(5'b00000),
	.iointdqslogicaclrpstamble(5'b00000),
	.iointdqslogicdqsena({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicfiforeset({gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincrdataen({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincwrptr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicoct({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicreadlatency({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointodtaclr(2'b00),
	.iointodtdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointrasndout({gnd,gnd,gnd,gnd}),
	.iointresetndout({gnd,gnd,gnd,gnd}),
	.iointwendout({gnd,gnd,gnd,gnd}),
	.aficalfail(afi_cal_fail),
	.aficalsuccess(afi_cal_success),
	.afirdatavalid(afi_rdata_valid[0]),
	.avlwaitrequest(),
	.ctlresetn(ctl_reset_n),
	.iointaficalfail(),
	.iointaficalsuccess(),
	.phyddiocasnaclr(),
	.phyddiorasnaclr(),
	.phyddioresetnaclr(),
	.phyddiowenaclr(),
	.phyresetn(),
	.afirdata(hphy_inst_AFIRDATA_bus),
	.afirlat(),
	.afiwlat(hphy_inst_AFIWLAT_bus),
	.avlreaddata(),
	.iointafirlat(),
	.iointafiwlat(),
	.iointdqdin(),
	.iointdqslogicrdatavalid(),
	.phyddioaddraclr(),
	.phyddioaddrdout(hphy_inst_PHYDDIOADDRDOUT_bus),
	.phyddiobaaclr(),
	.phyddiobadout(hphy_inst_PHYDDIOBADOUT_bus),
	.phyddiocasndout(hphy_inst_PHYDDIOCASNDOUT_bus),
	.phyddiockdout(hphy_inst_PHYDDIOCKDOUT_bus),
	.phyddiockeaclr(),
	.phyddiockedout(hphy_inst_PHYDDIOCKEDOUT_bus),
	.phyddiockndout(),
	.phyddiocsnaclr(),
	.phyddiocsndout(hphy_inst_PHYDDIOCSNDOUT_bus),
	.phyddiodmdout(hphy_inst_PHYDDIODMDOUT_bus),
	.phyddiodqdout(hphy_inst_PHYDDIODQDOUT_bus),
	.phyddiodqoe(hphy_inst_PHYDDIODQOE_bus),
	.phyddiodqsbdout(),
	.phyddiodqsboe(),
	.phyddiodqsdout(hphy_inst_PHYDDIODQSDOUT_bus),
	.phyddiodqslogicaclrfifoctrl(hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus),
	.phyddiodqslogicaclrpstamble(hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus),
	.phyddiodqslogicdqsena(hphy_inst_PHYDDIODQSLOGICDQSENA_bus),
	.phyddiodqslogicfiforeset(hphy_inst_PHYDDIODQSLOGICFIFORESET_bus),
	.phyddiodqslogicincrdataen(hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus),
	.phyddiodqslogicincwrptr(hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus),
	.phyddiodqslogicoct(hphy_inst_PHYDDIODQSLOGICOCT_bus),
	.phyddiodqslogicreadlatency(hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus),
	.phyddiodqsoe(hphy_inst_PHYDDIODQSOE_bus),
	.phyddioodtaclr(),
	.phyddioodtdout(hphy_inst_PHYDDIOODTDOUT_bus),
	.phyddiorasndout(hphy_inst_PHYDDIORASNDOUT_bus),
	.phyddioresetndout(hphy_inst_PHYDDIORESETNDOUT_bus),
	.phyddiowendout(hphy_inst_PHYDDIOWENDOUT_bus));
defparam hphy_inst.hphy_ac_ddr_disable = "true";
defparam hphy_inst.hphy_atpg_en = "false";
defparam hphy_inst.hphy_csr_pipelineglobalenable = "true";
defparam hphy_inst.hphy_datapath_ac_delay = "one_and_half_cycles";
defparam hphy_inst.hphy_datapath_delay = "one_cycle";
defparam hphy_inst.hphy_reset_delay_en = "false";
defparam hphy_inst.hphy_use_hphy = "true";
defparam hphy_inst.hphy_wrap_back_en = "false";
defparam hphy_inst.m_hphy_ac_rom_content = 1200'b100000011100000000000000000000100000011110000000000000000000010000000010000000010000110001010000000010000000010100110000010000000010010000000001000100010000000010100000000000010000010000000010110000000000000000010000001110000000010000000000010000000010000000010001001001010000000010000000010011001000010000000010100000000000100100010000000010010000000000001000010000000010110000000000000000110000011110000000000000000000111000011110000000000000000000110000011110000000000000000000010000011010000000000000000000010000011010110000000000000000010000001010000000010000000000010000010010000000000000000000011100100110000000000000000000011100100110110000000000000000011100100110000000000000001000011100100110110000000000001000111000111110000000000000000000111100111110000000000000000000111000011110000000000000000000011000000110000000000000000000011000100110000000000000000000010011010110000000000000000000010011010110110000000000000000010011010110000000000000001000010011010110110000000000001000110011011110000000000000000000010000010110000000000000001000010000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam hphy_inst.m_hphy_ac_rom_init_file = "hps_ac_rom.hex";
defparam hphy_inst.m_hphy_inst_rom_content = 2560'b1000000000000000000010000000011010000000000010000001100000000000100000100000000000001000001010000000000010000011000000000000100000111000000000001000000100000000000010000100100000000000100001010000000000001000010110000000000010000110000000000000100001000000000000000000100000000000000010000110100000000000000010001000000000001010011010000000100000000110100000000000000010010000000010000000011010000000000000001001100000000000101001101000000000001000011010000000100000000110100000000000000010110110100000001100110011101000000000001010111010000000100011001110100000000000101110001000000011101100100010000000000010100000100000001010110010001000100000000110100000000000110011100000000000001100110110000000000011100111000000000000000011000000000000100000110011100000001000001100111000000010000011001110000000100000110011100000000000001101000000000000000001101000000000000000011010000000000000000110100000000000000001101000000001100000111010000000011000010000100000000110000100001000000001100001000010000000000010100110100000000000100001101000000010000000011010000000000011001110000000000000110011011000000000001110011100000000000000001100000000000011000011001110000000110000110011100000001100001100111000000011000011001110000000000000110100000000000000000110100000000000000001101000000000000000011010000000000000000110100000000111000011101000000001110001000010000000011100010000100000000111000100001000000000001010011010000000000010000110100000001000000001101000000000000001000101011000000000000110110110001000000001101000000000000001000101101000000000000111111010000000000001111110100000001000011111101000010000001111111010000100000100001110100001000001000011101000010000010000111010000000000100010110100000000000011111101000000000000111111010000000101001111110100010000000011010000000010000001110100010000100000100001000100001000001000010001000010000010000100010000100000011110110100001000001000011101000010000010000111010000100000100001110100000001010011010000000010000001111111010000100000100001110100001000001000011101000010000010000111010000100000100000000100001000001000010001000010000010000100010000100000100001000100000000001000100000000000011000110100000000000100001101000000000001110011010000000100000000110100000000000000000000000000000001000000000000000000010100000000000000000110000000000000010000000000000000000000000000000100000000000100000001000000000001010000010000000000011000000100000001000000000001000000000001001000110000000000010000110100000000000101001101000000010000000011010000000010000001111000010001000000001101000000000000000000000000000;
defparam hphy_inst.m_hphy_inst_rom_init_file = "hps_inst_rom.hex";

endmodule

module soc_system_hps_sdram_p0_acv_hard_io_pads (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	input_path_gen0read_fifo_out_01,
	input_path_gen0read_fifo_out_11,
	input_path_gen0read_fifo_out_21,
	input_path_gen0read_fifo_out_31,
	input_path_gen1read_fifo_out_01,
	input_path_gen1read_fifo_out_11,
	input_path_gen1read_fifo_out_21,
	input_path_gen1read_fifo_out_31,
	input_path_gen2read_fifo_out_01,
	input_path_gen2read_fifo_out_11,
	input_path_gen2read_fifo_out_21,
	input_path_gen2read_fifo_out_31,
	input_path_gen3read_fifo_out_01,
	input_path_gen3read_fifo_out_11,
	input_path_gen3read_fifo_out_21,
	input_path_gen3read_fifo_out_31,
	input_path_gen4read_fifo_out_01,
	input_path_gen4read_fifo_out_11,
	input_path_gen4read_fifo_out_21,
	input_path_gen4read_fifo_out_31,
	input_path_gen5read_fifo_out_01,
	input_path_gen5read_fifo_out_11,
	input_path_gen5read_fifo_out_21,
	input_path_gen5read_fifo_out_31,
	input_path_gen6read_fifo_out_01,
	input_path_gen6read_fifo_out_11,
	input_path_gen6read_fifo_out_21,
	input_path_gen6read_fifo_out_31,
	input_path_gen7read_fifo_out_01,
	input_path_gen7read_fifo_out_11,
	input_path_gen7read_fifo_out_21,
	input_path_gen7read_fifo_out_31,
	input_path_gen0read_fifo_out_02,
	input_path_gen0read_fifo_out_12,
	input_path_gen0read_fifo_out_22,
	input_path_gen0read_fifo_out_32,
	input_path_gen1read_fifo_out_02,
	input_path_gen1read_fifo_out_12,
	input_path_gen1read_fifo_out_22,
	input_path_gen1read_fifo_out_32,
	input_path_gen2read_fifo_out_02,
	input_path_gen2read_fifo_out_12,
	input_path_gen2read_fifo_out_22,
	input_path_gen2read_fifo_out_32,
	input_path_gen3read_fifo_out_02,
	input_path_gen3read_fifo_out_12,
	input_path_gen3read_fifo_out_22,
	input_path_gen3read_fifo_out_32,
	input_path_gen4read_fifo_out_02,
	input_path_gen4read_fifo_out_12,
	input_path_gen4read_fifo_out_22,
	input_path_gen4read_fifo_out_32,
	input_path_gen5read_fifo_out_02,
	input_path_gen5read_fifo_out_12,
	input_path_gen5read_fifo_out_22,
	input_path_gen5read_fifo_out_32,
	input_path_gen6read_fifo_out_02,
	input_path_gen6read_fifo_out_12,
	input_path_gen6read_fifo_out_22,
	input_path_gen6read_fifo_out_32,
	input_path_gen7read_fifo_out_02,
	input_path_gen7read_fifo_out_12,
	input_path_gen7read_fifo_out_22,
	input_path_gen7read_fifo_out_32,
	input_path_gen0read_fifo_out_03,
	input_path_gen0read_fifo_out_13,
	input_path_gen0read_fifo_out_23,
	input_path_gen0read_fifo_out_33,
	input_path_gen1read_fifo_out_03,
	input_path_gen1read_fifo_out_13,
	input_path_gen1read_fifo_out_23,
	input_path_gen1read_fifo_out_33,
	input_path_gen2read_fifo_out_03,
	input_path_gen2read_fifo_out_13,
	input_path_gen2read_fifo_out_23,
	input_path_gen2read_fifo_out_33,
	input_path_gen3read_fifo_out_03,
	input_path_gen3read_fifo_out_13,
	input_path_gen3read_fifo_out_23,
	input_path_gen3read_fifo_out_33,
	input_path_gen4read_fifo_out_03,
	input_path_gen4read_fifo_out_13,
	input_path_gen4read_fifo_out_23,
	input_path_gen4read_fifo_out_33,
	input_path_gen5read_fifo_out_03,
	input_path_gen5read_fifo_out_13,
	input_path_gen5read_fifo_out_23,
	input_path_gen5read_fifo_out_33,
	input_path_gen6read_fifo_out_03,
	input_path_gen6read_fifo_out_13,
	input_path_gen6read_fifo_out_23,
	input_path_gen6read_fifo_out_33,
	input_path_gen7read_fifo_out_03,
	input_path_gen7read_fifo_out_13,
	input_path_gen7read_fifo_out_23,
	input_path_gen7read_fifo_out_33,
	ddio_phy_dqslogic_rdatavalid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	input_path_gen0read_fifo_out_01;
output 	input_path_gen0read_fifo_out_11;
output 	input_path_gen0read_fifo_out_21;
output 	input_path_gen0read_fifo_out_31;
output 	input_path_gen1read_fifo_out_01;
output 	input_path_gen1read_fifo_out_11;
output 	input_path_gen1read_fifo_out_21;
output 	input_path_gen1read_fifo_out_31;
output 	input_path_gen2read_fifo_out_01;
output 	input_path_gen2read_fifo_out_11;
output 	input_path_gen2read_fifo_out_21;
output 	input_path_gen2read_fifo_out_31;
output 	input_path_gen3read_fifo_out_01;
output 	input_path_gen3read_fifo_out_11;
output 	input_path_gen3read_fifo_out_21;
output 	input_path_gen3read_fifo_out_31;
output 	input_path_gen4read_fifo_out_01;
output 	input_path_gen4read_fifo_out_11;
output 	input_path_gen4read_fifo_out_21;
output 	input_path_gen4read_fifo_out_31;
output 	input_path_gen5read_fifo_out_01;
output 	input_path_gen5read_fifo_out_11;
output 	input_path_gen5read_fifo_out_21;
output 	input_path_gen5read_fifo_out_31;
output 	input_path_gen6read_fifo_out_01;
output 	input_path_gen6read_fifo_out_11;
output 	input_path_gen6read_fifo_out_21;
output 	input_path_gen6read_fifo_out_31;
output 	input_path_gen7read_fifo_out_01;
output 	input_path_gen7read_fifo_out_11;
output 	input_path_gen7read_fifo_out_21;
output 	input_path_gen7read_fifo_out_31;
output 	input_path_gen0read_fifo_out_02;
output 	input_path_gen0read_fifo_out_12;
output 	input_path_gen0read_fifo_out_22;
output 	input_path_gen0read_fifo_out_32;
output 	input_path_gen1read_fifo_out_02;
output 	input_path_gen1read_fifo_out_12;
output 	input_path_gen1read_fifo_out_22;
output 	input_path_gen1read_fifo_out_32;
output 	input_path_gen2read_fifo_out_02;
output 	input_path_gen2read_fifo_out_12;
output 	input_path_gen2read_fifo_out_22;
output 	input_path_gen2read_fifo_out_32;
output 	input_path_gen3read_fifo_out_02;
output 	input_path_gen3read_fifo_out_12;
output 	input_path_gen3read_fifo_out_22;
output 	input_path_gen3read_fifo_out_32;
output 	input_path_gen4read_fifo_out_02;
output 	input_path_gen4read_fifo_out_12;
output 	input_path_gen4read_fifo_out_22;
output 	input_path_gen4read_fifo_out_32;
output 	input_path_gen5read_fifo_out_02;
output 	input_path_gen5read_fifo_out_12;
output 	input_path_gen5read_fifo_out_22;
output 	input_path_gen5read_fifo_out_32;
output 	input_path_gen6read_fifo_out_02;
output 	input_path_gen6read_fifo_out_12;
output 	input_path_gen6read_fifo_out_22;
output 	input_path_gen6read_fifo_out_32;
output 	input_path_gen7read_fifo_out_02;
output 	input_path_gen7read_fifo_out_12;
output 	input_path_gen7read_fifo_out_22;
output 	input_path_gen7read_fifo_out_32;
output 	input_path_gen0read_fifo_out_03;
output 	input_path_gen0read_fifo_out_13;
output 	input_path_gen0read_fifo_out_23;
output 	input_path_gen0read_fifo_out_33;
output 	input_path_gen1read_fifo_out_03;
output 	input_path_gen1read_fifo_out_13;
output 	input_path_gen1read_fifo_out_23;
output 	input_path_gen1read_fifo_out_33;
output 	input_path_gen2read_fifo_out_03;
output 	input_path_gen2read_fifo_out_13;
output 	input_path_gen2read_fifo_out_23;
output 	input_path_gen2read_fifo_out_33;
output 	input_path_gen3read_fifo_out_03;
output 	input_path_gen3read_fifo_out_13;
output 	input_path_gen3read_fifo_out_23;
output 	input_path_gen3read_fifo_out_33;
output 	input_path_gen4read_fifo_out_03;
output 	input_path_gen4read_fifo_out_13;
output 	input_path_gen4read_fifo_out_23;
output 	input_path_gen4read_fifo_out_33;
output 	input_path_gen5read_fifo_out_03;
output 	input_path_gen5read_fifo_out_13;
output 	input_path_gen5read_fifo_out_23;
output 	input_path_gen5read_fifo_out_33;
output 	input_path_gen6read_fifo_out_03;
output 	input_path_gen6read_fifo_out_13;
output 	input_path_gen6read_fifo_out_23;
output 	input_path_gen6read_fifo_out_33;
output 	input_path_gen7read_fifo_out_03;
output 	input_path_gen7read_fifo_out_13;
output 	input_path_gen7read_fifo_out_23;
output 	input_path_gen7read_fifo_out_33;
output 	[4:0] ddio_phy_dqslogic_rdatavalid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_hps_sdram_p0_acv_hard_addr_cmd_pads uaddr_cmd_pads(
	.afi_clk(afi_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(phy_ddio_address_0),
	.phy_ddio_address_1(phy_ddio_address_1),
	.phy_ddio_address_2(phy_ddio_address_2),
	.phy_ddio_address_3(phy_ddio_address_3),
	.phy_ddio_address_4(phy_ddio_address_4),
	.phy_ddio_address_5(phy_ddio_address_5),
	.phy_ddio_address_6(phy_ddio_address_6),
	.phy_ddio_address_7(phy_ddio_address_7),
	.phy_ddio_address_8(phy_ddio_address_8),
	.phy_ddio_address_9(phy_ddio_address_9),
	.phy_ddio_address_10(phy_ddio_address_10),
	.phy_ddio_address_11(phy_ddio_address_11),
	.phy_ddio_address_12(phy_ddio_address_12),
	.phy_ddio_address_13(phy_ddio_address_13),
	.phy_ddio_address_14(phy_ddio_address_14),
	.phy_ddio_address_15(phy_ddio_address_15),
	.phy_ddio_address_16(phy_ddio_address_16),
	.phy_ddio_address_17(phy_ddio_address_17),
	.phy_ddio_address_18(phy_ddio_address_18),
	.phy_ddio_address_19(phy_ddio_address_19),
	.phy_ddio_address_20(phy_ddio_address_20),
	.phy_ddio_address_21(phy_ddio_address_21),
	.phy_ddio_address_22(phy_ddio_address_22),
	.phy_ddio_address_23(phy_ddio_address_23),
	.phy_ddio_address_24(phy_ddio_address_24),
	.phy_ddio_address_25(phy_ddio_address_25),
	.phy_ddio_address_26(phy_ddio_address_26),
	.phy_ddio_address_27(phy_ddio_address_27),
	.phy_ddio_address_28(phy_ddio_address_28),
	.phy_ddio_address_29(phy_ddio_address_29),
	.phy_ddio_address_30(phy_ddio_address_30),
	.phy_ddio_address_31(phy_ddio_address_31),
	.phy_ddio_address_32(phy_ddio_address_32),
	.phy_ddio_address_33(phy_ddio_address_33),
	.phy_ddio_address_34(phy_ddio_address_34),
	.phy_ddio_address_35(phy_ddio_address_35),
	.phy_ddio_address_36(phy_ddio_address_36),
	.phy_ddio_address_37(phy_ddio_address_37),
	.phy_ddio_address_38(phy_ddio_address_38),
	.phy_ddio_address_39(phy_ddio_address_39),
	.phy_ddio_address_40(phy_ddio_address_40),
	.phy_ddio_address_41(phy_ddio_address_41),
	.phy_ddio_address_42(phy_ddio_address_42),
	.phy_ddio_address_43(phy_ddio_address_43),
	.phy_ddio_address_44(phy_ddio_address_44),
	.phy_ddio_address_45(phy_ddio_address_45),
	.phy_ddio_address_46(phy_ddio_address_46),
	.phy_ddio_address_47(phy_ddio_address_47),
	.phy_ddio_address_48(phy_ddio_address_48),
	.phy_ddio_address_49(phy_ddio_address_49),
	.phy_ddio_address_50(phy_ddio_address_50),
	.phy_ddio_address_51(phy_ddio_address_51),
	.phy_ddio_address_52(phy_ddio_address_52),
	.phy_ddio_address_53(phy_ddio_address_53),
	.phy_ddio_address_54(phy_ddio_address_54),
	.phy_ddio_address_55(phy_ddio_address_55),
	.phy_ddio_address_56(phy_ddio_address_56),
	.phy_ddio_address_57(phy_ddio_address_57),
	.phy_ddio_address_58(phy_ddio_address_58),
	.phy_ddio_address_59(phy_ddio_address_59),
	.phy_ddio_bank_0(phy_ddio_bank_0),
	.phy_ddio_bank_1(phy_ddio_bank_1),
	.phy_ddio_bank_2(phy_ddio_bank_2),
	.phy_ddio_bank_3(phy_ddio_bank_3),
	.phy_ddio_bank_4(phy_ddio_bank_4),
	.phy_ddio_bank_5(phy_ddio_bank_5),
	.phy_ddio_bank_6(phy_ddio_bank_6),
	.phy_ddio_bank_7(phy_ddio_bank_7),
	.phy_ddio_bank_8(phy_ddio_bank_8),
	.phy_ddio_bank_9(phy_ddio_bank_9),
	.phy_ddio_bank_10(phy_ddio_bank_10),
	.phy_ddio_bank_11(phy_ddio_bank_11),
	.phy_ddio_cas_n_0(phy_ddio_cas_n_0),
	.phy_ddio_cas_n_1(phy_ddio_cas_n_1),
	.phy_ddio_cas_n_2(phy_ddio_cas_n_2),
	.phy_ddio_cas_n_3(phy_ddio_cas_n_3),
	.phy_ddio_ck_0(phy_ddio_ck_0),
	.phy_ddio_ck_1(phy_ddio_ck_1),
	.phy_ddio_cke_0(phy_ddio_cke_0),
	.phy_ddio_cke_1(phy_ddio_cke_1),
	.phy_ddio_cke_2(phy_ddio_cke_2),
	.phy_ddio_cke_3(phy_ddio_cke_3),
	.phy_ddio_cs_n_0(phy_ddio_cs_n_0),
	.phy_ddio_cs_n_1(phy_ddio_cs_n_1),
	.phy_ddio_cs_n_2(phy_ddio_cs_n_2),
	.phy_ddio_cs_n_3(phy_ddio_cs_n_3),
	.phy_ddio_odt_0(phy_ddio_odt_0),
	.phy_ddio_odt_1(phy_ddio_odt_1),
	.phy_ddio_odt_2(phy_ddio_odt_2),
	.phy_ddio_odt_3(phy_ddio_odt_3),
	.phy_ddio_ras_n_0(phy_ddio_ras_n_0),
	.phy_ddio_ras_n_1(phy_ddio_ras_n_1),
	.phy_ddio_ras_n_2(phy_ddio_ras_n_2),
	.phy_ddio_ras_n_3(phy_ddio_ras_n_3),
	.phy_ddio_reset_n_0(phy_ddio_reset_n_0),
	.phy_ddio_reset_n_1(phy_ddio_reset_n_1),
	.phy_ddio_reset_n_2(phy_ddio_reset_n_2),
	.phy_ddio_reset_n_3(phy_ddio_reset_n_3),
	.phy_ddio_we_n_0(phy_ddio_we_n_0),
	.phy_ddio_we_n_1(phy_ddio_we_n_1),
	.phy_ddio_we_n_2(phy_ddio_we_n_2),
	.phy_ddio_we_n_3(phy_ddio_we_n_3),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6));

soc_system_hps_sdram_p0_altdqdqs_3 \dq_ddio[3].ubidir_dq_dqs (
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.phy_ddio_dmdout_12(phy_ddio_dmdout_12),
	.phy_ddio_dmdout_13(phy_ddio_dmdout_13),
	.phy_ddio_dmdout_14(phy_ddio_dmdout_14),
	.phy_ddio_dmdout_15(phy_ddio_dmdout_15),
	.phy_ddio_dqdout_108(phy_ddio_dqdout_108),
	.phy_ddio_dqdout_109(phy_ddio_dqdout_109),
	.phy_ddio_dqdout_110(phy_ddio_dqdout_110),
	.phy_ddio_dqdout_111(phy_ddio_dqdout_111),
	.phy_ddio_dqdout_112(phy_ddio_dqdout_112),
	.phy_ddio_dqdout_113(phy_ddio_dqdout_113),
	.phy_ddio_dqdout_114(phy_ddio_dqdout_114),
	.phy_ddio_dqdout_115(phy_ddio_dqdout_115),
	.phy_ddio_dqdout_116(phy_ddio_dqdout_116),
	.phy_ddio_dqdout_117(phy_ddio_dqdout_117),
	.phy_ddio_dqdout_118(phy_ddio_dqdout_118),
	.phy_ddio_dqdout_119(phy_ddio_dqdout_119),
	.phy_ddio_dqdout_120(phy_ddio_dqdout_120),
	.phy_ddio_dqdout_121(phy_ddio_dqdout_121),
	.phy_ddio_dqdout_122(phy_ddio_dqdout_122),
	.phy_ddio_dqdout_123(phy_ddio_dqdout_123),
	.phy_ddio_dqdout_124(phy_ddio_dqdout_124),
	.phy_ddio_dqdout_125(phy_ddio_dqdout_125),
	.phy_ddio_dqdout_126(phy_ddio_dqdout_126),
	.phy_ddio_dqdout_127(phy_ddio_dqdout_127),
	.phy_ddio_dqdout_128(phy_ddio_dqdout_128),
	.phy_ddio_dqdout_129(phy_ddio_dqdout_129),
	.phy_ddio_dqdout_130(phy_ddio_dqdout_130),
	.phy_ddio_dqdout_131(phy_ddio_dqdout_131),
	.phy_ddio_dqdout_132(phy_ddio_dqdout_132),
	.phy_ddio_dqdout_133(phy_ddio_dqdout_133),
	.phy_ddio_dqdout_134(phy_ddio_dqdout_134),
	.phy_ddio_dqdout_135(phy_ddio_dqdout_135),
	.phy_ddio_dqdout_136(phy_ddio_dqdout_136),
	.phy_ddio_dqdout_137(phy_ddio_dqdout_137),
	.phy_ddio_dqdout_138(phy_ddio_dqdout_138),
	.phy_ddio_dqdout_139(phy_ddio_dqdout_139),
	.phy_ddio_dqoe_54(phy_ddio_dqoe_54),
	.phy_ddio_dqoe_55(phy_ddio_dqoe_55),
	.phy_ddio_dqoe_56(phy_ddio_dqoe_56),
	.phy_ddio_dqoe_57(phy_ddio_dqoe_57),
	.phy_ddio_dqoe_58(phy_ddio_dqoe_58),
	.phy_ddio_dqoe_59(phy_ddio_dqoe_59),
	.phy_ddio_dqoe_60(phy_ddio_dqoe_60),
	.phy_ddio_dqoe_61(phy_ddio_dqoe_61),
	.phy_ddio_dqoe_62(phy_ddio_dqoe_62),
	.phy_ddio_dqoe_63(phy_ddio_dqoe_63),
	.phy_ddio_dqoe_64(phy_ddio_dqoe_64),
	.phy_ddio_dqoe_65(phy_ddio_dqoe_65),
	.phy_ddio_dqoe_66(phy_ddio_dqoe_66),
	.phy_ddio_dqoe_67(phy_ddio_dqoe_67),
	.phy_ddio_dqoe_68(phy_ddio_dqoe_68),
	.phy_ddio_dqoe_69(phy_ddio_dqoe_69),
	.phy_ddio_dqs_dout_12(phy_ddio_dqs_dout_12),
	.phy_ddio_dqs_dout_13(phy_ddio_dqs_dout_13),
	.phy_ddio_dqs_dout_14(phy_ddio_dqs_dout_14),
	.phy_ddio_dqs_dout_15(phy_ddio_dqs_dout_15),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.phy_ddio_dqslogic_aclr_pstamble_3(phy_ddio_dqslogic_aclr_pstamble_3),
	.phy_ddio_dqslogic_dqsena_6(phy_ddio_dqslogic_dqsena_6),
	.phy_ddio_dqslogic_dqsena_7(phy_ddio_dqslogic_dqsena_7),
	.phy_ddio_dqslogic_fiforeset_3(phy_ddio_dqslogic_fiforeset_3),
	.phy_ddio_dqslogic_incrdataen_6(phy_ddio_dqslogic_incrdataen_6),
	.phy_ddio_dqslogic_incrdataen_7(phy_ddio_dqslogic_incrdataen_7),
	.phy_ddio_dqslogic_incwrptr_6(phy_ddio_dqslogic_incwrptr_6),
	.phy_ddio_dqslogic_incwrptr_7(phy_ddio_dqslogic_incwrptr_7),
	.phy_ddio_dqslogic_oct_6(phy_ddio_dqslogic_oct_6),
	.phy_ddio_dqslogic_oct_7(phy_ddio_dqslogic_oct_7),
	.phy_ddio_dqslogic_readlatency_15(phy_ddio_dqslogic_readlatency_15),
	.phy_ddio_dqslogic_readlatency_16(phy_ddio_dqslogic_readlatency_16),
	.phy_ddio_dqslogic_readlatency_17(phy_ddio_dqslogic_readlatency_17),
	.phy_ddio_dqslogic_readlatency_18(phy_ddio_dqslogic_readlatency_18),
	.phy_ddio_dqslogic_readlatency_19(phy_ddio_dqslogic_readlatency_19),
	.phy_ddio_dqs_oe_6(phy_ddio_dqs_oe_6),
	.phy_ddio_dqs_oe_7(phy_ddio_dqs_oe_7),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_13),
	.delayed_oct(delayed_oct3),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_13),
	.os(os3),
	.os_bar(os_bar3),
	.diff_oe(diff_oe3),
	.diff_oe_bar(diff_oe_bar3),
	.diff_dtc(diff_dtc3),
	.diff_dtc_bar(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_03),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_13),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_23),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_33),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_03),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_13),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_23),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_33),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_03),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_13),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_23),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_33),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_03),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_13),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_23),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_33),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_03),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_13),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_23),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_33),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_03),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_13),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_23),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_33),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_03),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_13),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_23),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_33),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_03),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_13),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_23),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_33),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[3]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

soc_system_hps_sdram_p0_altdqdqs_2 \dq_ddio[2].ubidir_dq_dqs (
	.dqsin(dqsin1),
	.pad_gen0raw_input(pad_gen0raw_input1),
	.pad_gen1raw_input(pad_gen1raw_input1),
	.pad_gen2raw_input(pad_gen2raw_input1),
	.pad_gen3raw_input(pad_gen3raw_input1),
	.pad_gen4raw_input(pad_gen4raw_input1),
	.pad_gen5raw_input(pad_gen5raw_input1),
	.pad_gen6raw_input(pad_gen6raw_input1),
	.pad_gen7raw_input(pad_gen7raw_input1),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out1),
	.phy_ddio_dmdout_8(phy_ddio_dmdout_8),
	.phy_ddio_dmdout_9(phy_ddio_dmdout_9),
	.phy_ddio_dmdout_10(phy_ddio_dmdout_10),
	.phy_ddio_dmdout_11(phy_ddio_dmdout_11),
	.phy_ddio_dqdout_72(phy_ddio_dqdout_72),
	.phy_ddio_dqdout_73(phy_ddio_dqdout_73),
	.phy_ddio_dqdout_74(phy_ddio_dqdout_74),
	.phy_ddio_dqdout_75(phy_ddio_dqdout_75),
	.phy_ddio_dqdout_76(phy_ddio_dqdout_76),
	.phy_ddio_dqdout_77(phy_ddio_dqdout_77),
	.phy_ddio_dqdout_78(phy_ddio_dqdout_78),
	.phy_ddio_dqdout_79(phy_ddio_dqdout_79),
	.phy_ddio_dqdout_80(phy_ddio_dqdout_80),
	.phy_ddio_dqdout_81(phy_ddio_dqdout_81),
	.phy_ddio_dqdout_82(phy_ddio_dqdout_82),
	.phy_ddio_dqdout_83(phy_ddio_dqdout_83),
	.phy_ddio_dqdout_84(phy_ddio_dqdout_84),
	.phy_ddio_dqdout_85(phy_ddio_dqdout_85),
	.phy_ddio_dqdout_86(phy_ddio_dqdout_86),
	.phy_ddio_dqdout_87(phy_ddio_dqdout_87),
	.phy_ddio_dqdout_88(phy_ddio_dqdout_88),
	.phy_ddio_dqdout_89(phy_ddio_dqdout_89),
	.phy_ddio_dqdout_90(phy_ddio_dqdout_90),
	.phy_ddio_dqdout_91(phy_ddio_dqdout_91),
	.phy_ddio_dqdout_92(phy_ddio_dqdout_92),
	.phy_ddio_dqdout_93(phy_ddio_dqdout_93),
	.phy_ddio_dqdout_94(phy_ddio_dqdout_94),
	.phy_ddio_dqdout_95(phy_ddio_dqdout_95),
	.phy_ddio_dqdout_96(phy_ddio_dqdout_96),
	.phy_ddio_dqdout_97(phy_ddio_dqdout_97),
	.phy_ddio_dqdout_98(phy_ddio_dqdout_98),
	.phy_ddio_dqdout_99(phy_ddio_dqdout_99),
	.phy_ddio_dqdout_100(phy_ddio_dqdout_100),
	.phy_ddio_dqdout_101(phy_ddio_dqdout_101),
	.phy_ddio_dqdout_102(phy_ddio_dqdout_102),
	.phy_ddio_dqdout_103(phy_ddio_dqdout_103),
	.phy_ddio_dqoe_36(phy_ddio_dqoe_36),
	.phy_ddio_dqoe_37(phy_ddio_dqoe_37),
	.phy_ddio_dqoe_38(phy_ddio_dqoe_38),
	.phy_ddio_dqoe_39(phy_ddio_dqoe_39),
	.phy_ddio_dqoe_40(phy_ddio_dqoe_40),
	.phy_ddio_dqoe_41(phy_ddio_dqoe_41),
	.phy_ddio_dqoe_42(phy_ddio_dqoe_42),
	.phy_ddio_dqoe_43(phy_ddio_dqoe_43),
	.phy_ddio_dqoe_44(phy_ddio_dqoe_44),
	.phy_ddio_dqoe_45(phy_ddio_dqoe_45),
	.phy_ddio_dqoe_46(phy_ddio_dqoe_46),
	.phy_ddio_dqoe_47(phy_ddio_dqoe_47),
	.phy_ddio_dqoe_48(phy_ddio_dqoe_48),
	.phy_ddio_dqoe_49(phy_ddio_dqoe_49),
	.phy_ddio_dqoe_50(phy_ddio_dqoe_50),
	.phy_ddio_dqoe_51(phy_ddio_dqoe_51),
	.phy_ddio_dqs_dout_8(phy_ddio_dqs_dout_8),
	.phy_ddio_dqs_dout_9(phy_ddio_dqs_dout_9),
	.phy_ddio_dqs_dout_10(phy_ddio_dqs_dout_10),
	.phy_ddio_dqs_dout_11(phy_ddio_dqs_dout_11),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.phy_ddio_dqslogic_aclr_pstamble_2(phy_ddio_dqslogic_aclr_pstamble_2),
	.phy_ddio_dqslogic_dqsena_4(phy_ddio_dqslogic_dqsena_4),
	.phy_ddio_dqslogic_dqsena_5(phy_ddio_dqslogic_dqsena_5),
	.phy_ddio_dqslogic_fiforeset_2(phy_ddio_dqslogic_fiforeset_2),
	.phy_ddio_dqslogic_incrdataen_4(phy_ddio_dqslogic_incrdataen_4),
	.phy_ddio_dqslogic_incrdataen_5(phy_ddio_dqslogic_incrdataen_5),
	.phy_ddio_dqslogic_incwrptr_4(phy_ddio_dqslogic_incwrptr_4),
	.phy_ddio_dqslogic_incwrptr_5(phy_ddio_dqslogic_incwrptr_5),
	.phy_ddio_dqslogic_oct_4(phy_ddio_dqslogic_oct_4),
	.phy_ddio_dqslogic_oct_5(phy_ddio_dqslogic_oct_5),
	.phy_ddio_dqslogic_readlatency_10(phy_ddio_dqslogic_readlatency_10),
	.phy_ddio_dqslogic_readlatency_11(phy_ddio_dqslogic_readlatency_11),
	.phy_ddio_dqslogic_readlatency_12(phy_ddio_dqslogic_readlatency_12),
	.phy_ddio_dqslogic_readlatency_13(phy_ddio_dqslogic_readlatency_13),
	.phy_ddio_dqslogic_readlatency_14(phy_ddio_dqslogic_readlatency_14),
	.phy_ddio_dqs_oe_4(phy_ddio_dqs_oe_4),
	.phy_ddio_dqs_oe_5(phy_ddio_dqs_oe_5),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_12),
	.delayed_oct(delayed_oct2),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_12),
	.os(os2),
	.os_bar(os_bar2),
	.diff_oe(diff_oe2),
	.diff_oe_bar(diff_oe_bar2),
	.diff_dtc(diff_dtc2),
	.diff_dtc_bar(diff_dtc_bar2),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_02),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_12),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_22),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_32),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_02),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_12),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_22),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_32),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_02),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_12),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_22),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_32),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_02),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_12),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_22),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_32),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_02),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_12),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_22),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_32),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_02),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_12),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_22),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_32),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_02),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_12),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_22),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_32),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_02),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_12),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_22),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_32),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[2]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

soc_system_hps_sdram_p0_altdqdqs_1 \dq_ddio[1].ubidir_dq_dqs (
	.dqsin(dqsin2),
	.pad_gen0raw_input(pad_gen0raw_input2),
	.pad_gen1raw_input(pad_gen1raw_input2),
	.pad_gen2raw_input(pad_gen2raw_input2),
	.pad_gen3raw_input(pad_gen3raw_input2),
	.pad_gen4raw_input(pad_gen4raw_input2),
	.pad_gen5raw_input(pad_gen5raw_input2),
	.pad_gen6raw_input(pad_gen6raw_input2),
	.pad_gen7raw_input(pad_gen7raw_input2),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out2),
	.phy_ddio_dmdout_4(phy_ddio_dmdout_4),
	.phy_ddio_dmdout_5(phy_ddio_dmdout_5),
	.phy_ddio_dmdout_6(phy_ddio_dmdout_6),
	.phy_ddio_dmdout_7(phy_ddio_dmdout_7),
	.phy_ddio_dqdout_36(phy_ddio_dqdout_36),
	.phy_ddio_dqdout_37(phy_ddio_dqdout_37),
	.phy_ddio_dqdout_38(phy_ddio_dqdout_38),
	.phy_ddio_dqdout_39(phy_ddio_dqdout_39),
	.phy_ddio_dqdout_40(phy_ddio_dqdout_40),
	.phy_ddio_dqdout_41(phy_ddio_dqdout_41),
	.phy_ddio_dqdout_42(phy_ddio_dqdout_42),
	.phy_ddio_dqdout_43(phy_ddio_dqdout_43),
	.phy_ddio_dqdout_44(phy_ddio_dqdout_44),
	.phy_ddio_dqdout_45(phy_ddio_dqdout_45),
	.phy_ddio_dqdout_46(phy_ddio_dqdout_46),
	.phy_ddio_dqdout_47(phy_ddio_dqdout_47),
	.phy_ddio_dqdout_48(phy_ddio_dqdout_48),
	.phy_ddio_dqdout_49(phy_ddio_dqdout_49),
	.phy_ddio_dqdout_50(phy_ddio_dqdout_50),
	.phy_ddio_dqdout_51(phy_ddio_dqdout_51),
	.phy_ddio_dqdout_52(phy_ddio_dqdout_52),
	.phy_ddio_dqdout_53(phy_ddio_dqdout_53),
	.phy_ddio_dqdout_54(phy_ddio_dqdout_54),
	.phy_ddio_dqdout_55(phy_ddio_dqdout_55),
	.phy_ddio_dqdout_56(phy_ddio_dqdout_56),
	.phy_ddio_dqdout_57(phy_ddio_dqdout_57),
	.phy_ddio_dqdout_58(phy_ddio_dqdout_58),
	.phy_ddio_dqdout_59(phy_ddio_dqdout_59),
	.phy_ddio_dqdout_60(phy_ddio_dqdout_60),
	.phy_ddio_dqdout_61(phy_ddio_dqdout_61),
	.phy_ddio_dqdout_62(phy_ddio_dqdout_62),
	.phy_ddio_dqdout_63(phy_ddio_dqdout_63),
	.phy_ddio_dqdout_64(phy_ddio_dqdout_64),
	.phy_ddio_dqdout_65(phy_ddio_dqdout_65),
	.phy_ddio_dqdout_66(phy_ddio_dqdout_66),
	.phy_ddio_dqdout_67(phy_ddio_dqdout_67),
	.phy_ddio_dqoe_18(phy_ddio_dqoe_18),
	.phy_ddio_dqoe_19(phy_ddio_dqoe_19),
	.phy_ddio_dqoe_20(phy_ddio_dqoe_20),
	.phy_ddio_dqoe_21(phy_ddio_dqoe_21),
	.phy_ddio_dqoe_22(phy_ddio_dqoe_22),
	.phy_ddio_dqoe_23(phy_ddio_dqoe_23),
	.phy_ddio_dqoe_24(phy_ddio_dqoe_24),
	.phy_ddio_dqoe_25(phy_ddio_dqoe_25),
	.phy_ddio_dqoe_26(phy_ddio_dqoe_26),
	.phy_ddio_dqoe_27(phy_ddio_dqoe_27),
	.phy_ddio_dqoe_28(phy_ddio_dqoe_28),
	.phy_ddio_dqoe_29(phy_ddio_dqoe_29),
	.phy_ddio_dqoe_30(phy_ddio_dqoe_30),
	.phy_ddio_dqoe_31(phy_ddio_dqoe_31),
	.phy_ddio_dqoe_32(phy_ddio_dqoe_32),
	.phy_ddio_dqoe_33(phy_ddio_dqoe_33),
	.phy_ddio_dqs_dout_4(phy_ddio_dqs_dout_4),
	.phy_ddio_dqs_dout_5(phy_ddio_dqs_dout_5),
	.phy_ddio_dqs_dout_6(phy_ddio_dqs_dout_6),
	.phy_ddio_dqs_dout_7(phy_ddio_dqs_dout_7),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.phy_ddio_dqslogic_aclr_pstamble_1(phy_ddio_dqslogic_aclr_pstamble_1),
	.phy_ddio_dqslogic_dqsena_2(phy_ddio_dqslogic_dqsena_2),
	.phy_ddio_dqslogic_dqsena_3(phy_ddio_dqslogic_dqsena_3),
	.phy_ddio_dqslogic_fiforeset_1(phy_ddio_dqslogic_fiforeset_1),
	.phy_ddio_dqslogic_incrdataen_2(phy_ddio_dqslogic_incrdataen_2),
	.phy_ddio_dqslogic_incrdataen_3(phy_ddio_dqslogic_incrdataen_3),
	.phy_ddio_dqslogic_incwrptr_2(phy_ddio_dqslogic_incwrptr_2),
	.phy_ddio_dqslogic_incwrptr_3(phy_ddio_dqslogic_incwrptr_3),
	.phy_ddio_dqslogic_oct_2(phy_ddio_dqslogic_oct_2),
	.phy_ddio_dqslogic_oct_3(phy_ddio_dqslogic_oct_3),
	.phy_ddio_dqslogic_readlatency_5(phy_ddio_dqslogic_readlatency_5),
	.phy_ddio_dqslogic_readlatency_6(phy_ddio_dqslogic_readlatency_6),
	.phy_ddio_dqslogic_readlatency_7(phy_ddio_dqslogic_readlatency_7),
	.phy_ddio_dqslogic_readlatency_8(phy_ddio_dqslogic_readlatency_8),
	.phy_ddio_dqslogic_readlatency_9(phy_ddio_dqslogic_readlatency_9),
	.phy_ddio_dqs_oe_2(phy_ddio_dqs_oe_2),
	.phy_ddio_dqs_oe_3(phy_ddio_dqs_oe_3),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_11),
	.delayed_oct(delayed_oct1),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_11),
	.os(os1),
	.os_bar(os_bar1),
	.diff_oe(diff_oe1),
	.diff_oe_bar(diff_oe_bar1),
	.diff_dtc(diff_dtc1),
	.diff_dtc_bar(diff_dtc_bar1),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_01),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_11),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_21),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_31),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_01),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_11),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_21),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_31),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_01),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_11),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_21),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_31),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_01),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_11),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_21),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_31),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_01),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_11),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_21),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_31),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_01),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_11),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_21),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_31),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_01),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_11),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_21),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_31),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_01),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_11),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_21),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_31),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[1]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

soc_system_hps_sdram_p0_altdqdqs \dq_ddio[0].ubidir_dq_dqs (
	.dqsin(dqsin3),
	.pad_gen0raw_input(pad_gen0raw_input3),
	.pad_gen1raw_input(pad_gen1raw_input3),
	.pad_gen2raw_input(pad_gen2raw_input3),
	.pad_gen3raw_input(pad_gen3raw_input3),
	.pad_gen4raw_input(pad_gen4raw_input3),
	.pad_gen5raw_input(pad_gen5raw_input3),
	.pad_gen6raw_input(pad_gen6raw_input3),
	.pad_gen7raw_input(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out3),
	.phy_ddio_dmdout_0(phy_ddio_dmdout_0),
	.phy_ddio_dmdout_1(phy_ddio_dmdout_1),
	.phy_ddio_dmdout_2(phy_ddio_dmdout_2),
	.phy_ddio_dmdout_3(phy_ddio_dmdout_3),
	.phy_ddio_dqdout_0(phy_ddio_dqdout_0),
	.phy_ddio_dqdout_1(phy_ddio_dqdout_1),
	.phy_ddio_dqdout_2(phy_ddio_dqdout_2),
	.phy_ddio_dqdout_3(phy_ddio_dqdout_3),
	.phy_ddio_dqdout_4(phy_ddio_dqdout_4),
	.phy_ddio_dqdout_5(phy_ddio_dqdout_5),
	.phy_ddio_dqdout_6(phy_ddio_dqdout_6),
	.phy_ddio_dqdout_7(phy_ddio_dqdout_7),
	.phy_ddio_dqdout_8(phy_ddio_dqdout_8),
	.phy_ddio_dqdout_9(phy_ddio_dqdout_9),
	.phy_ddio_dqdout_10(phy_ddio_dqdout_10),
	.phy_ddio_dqdout_11(phy_ddio_dqdout_11),
	.phy_ddio_dqdout_12(phy_ddio_dqdout_12),
	.phy_ddio_dqdout_13(phy_ddio_dqdout_13),
	.phy_ddio_dqdout_14(phy_ddio_dqdout_14),
	.phy_ddio_dqdout_15(phy_ddio_dqdout_15),
	.phy_ddio_dqdout_16(phy_ddio_dqdout_16),
	.phy_ddio_dqdout_17(phy_ddio_dqdout_17),
	.phy_ddio_dqdout_18(phy_ddio_dqdout_18),
	.phy_ddio_dqdout_19(phy_ddio_dqdout_19),
	.phy_ddio_dqdout_20(phy_ddio_dqdout_20),
	.phy_ddio_dqdout_21(phy_ddio_dqdout_21),
	.phy_ddio_dqdout_22(phy_ddio_dqdout_22),
	.phy_ddio_dqdout_23(phy_ddio_dqdout_23),
	.phy_ddio_dqdout_24(phy_ddio_dqdout_24),
	.phy_ddio_dqdout_25(phy_ddio_dqdout_25),
	.phy_ddio_dqdout_26(phy_ddio_dqdout_26),
	.phy_ddio_dqdout_27(phy_ddio_dqdout_27),
	.phy_ddio_dqdout_28(phy_ddio_dqdout_28),
	.phy_ddio_dqdout_29(phy_ddio_dqdout_29),
	.phy_ddio_dqdout_30(phy_ddio_dqdout_30),
	.phy_ddio_dqdout_31(phy_ddio_dqdout_31),
	.phy_ddio_dqoe_0(phy_ddio_dqoe_0),
	.phy_ddio_dqoe_1(phy_ddio_dqoe_1),
	.phy_ddio_dqoe_2(phy_ddio_dqoe_2),
	.phy_ddio_dqoe_3(phy_ddio_dqoe_3),
	.phy_ddio_dqoe_4(phy_ddio_dqoe_4),
	.phy_ddio_dqoe_5(phy_ddio_dqoe_5),
	.phy_ddio_dqoe_6(phy_ddio_dqoe_6),
	.phy_ddio_dqoe_7(phy_ddio_dqoe_7),
	.phy_ddio_dqoe_8(phy_ddio_dqoe_8),
	.phy_ddio_dqoe_9(phy_ddio_dqoe_9),
	.phy_ddio_dqoe_10(phy_ddio_dqoe_10),
	.phy_ddio_dqoe_11(phy_ddio_dqoe_11),
	.phy_ddio_dqoe_12(phy_ddio_dqoe_12),
	.phy_ddio_dqoe_13(phy_ddio_dqoe_13),
	.phy_ddio_dqoe_14(phy_ddio_dqoe_14),
	.phy_ddio_dqoe_15(phy_ddio_dqoe_15),
	.phy_ddio_dqs_dout_0(phy_ddio_dqs_dout_0),
	.phy_ddio_dqs_dout_1(phy_ddio_dqs_dout_1),
	.phy_ddio_dqs_dout_2(phy_ddio_dqs_dout_2),
	.phy_ddio_dqs_dout_3(phy_ddio_dqs_dout_3),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.phy_ddio_dqslogic_aclr_pstamble_0(phy_ddio_dqslogic_aclr_pstamble_0),
	.phy_ddio_dqslogic_dqsena_0(phy_ddio_dqslogic_dqsena_0),
	.phy_ddio_dqslogic_dqsena_1(phy_ddio_dqslogic_dqsena_1),
	.phy_ddio_dqslogic_fiforeset_0(phy_ddio_dqslogic_fiforeset_0),
	.phy_ddio_dqslogic_incrdataen_0(phy_ddio_dqslogic_incrdataen_0),
	.phy_ddio_dqslogic_incrdataen_1(phy_ddio_dqslogic_incrdataen_1),
	.phy_ddio_dqslogic_incwrptr_0(phy_ddio_dqslogic_incwrptr_0),
	.phy_ddio_dqslogic_incwrptr_1(phy_ddio_dqslogic_incwrptr_1),
	.phy_ddio_dqslogic_oct_0(phy_ddio_dqslogic_oct_0),
	.phy_ddio_dqslogic_oct_1(phy_ddio_dqslogic_oct_1),
	.phy_ddio_dqslogic_readlatency_0(phy_ddio_dqslogic_readlatency_0),
	.phy_ddio_dqslogic_readlatency_1(phy_ddio_dqslogic_readlatency_1),
	.phy_ddio_dqslogic_readlatency_2(phy_ddio_dqslogic_readlatency_2),
	.phy_ddio_dqslogic_readlatency_3(phy_ddio_dqslogic_readlatency_3),
	.phy_ddio_dqslogic_readlatency_4(phy_ddio_dqslogic_readlatency_4),
	.phy_ddio_dqs_oe_0(phy_ddio_dqs_oe_0),
	.phy_ddio_dqs_oe_1(phy_ddio_dqs_oe_1),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_0),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_1),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_2),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_3),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_0),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_1),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_2),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_3),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_0),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_1),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_2),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_3),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_0),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_1),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_2),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_3),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_0),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_1),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_2),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_3),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_0),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_1),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_2),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_3),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_0),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_1),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_2),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_3),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_0),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_1),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_2),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_3),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[0]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module soc_system_hps_sdram_p0_acv_hard_addr_cmd_pads (
	afi_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6)/* synthesis synthesis_greybox=0 */;
input 	afi_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_gen[0].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[1].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[2].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[3].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[4].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[5].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[6].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[7].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[8].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[9].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[10].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[11].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[12].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[13].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[14].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[15].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[16].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[17].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[19].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[18].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[21].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[22].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[23].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[24].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[20].acv_ac_ldc|adc_clk_cps ;
wire \clock_gen[0].umem_ck_pad|auto_generated|dataout[0] ;
wire \mem_ck_source[0] ;
wire \clock_gen[0].leveled_dqs_clocks[0] ;
wire \clock_gen[0].leveled_dqs_clocks[1] ;
wire \clock_gen[0].leveled_dqs_clocks[2] ;
wire \clock_gen[0].leveled_dqs_clocks[3] ;

wire [3:0] \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ;

assign \clock_gen[0].leveled_dqs_clocks[0]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [0];
assign \clock_gen[0].leveled_dqs_clocks[1]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [1];
assign \clock_gen[0].leveled_dqs_clocks[2]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [2];
assign \clock_gen[0].leveled_dqs_clocks[3]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [3];

soc_system_hps_sdram_p0_acv_ldc_18 \address_gen[3].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[3].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_17 \address_gen[2].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[2].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_11 \address_gen[1].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[1].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc \address_gen[0].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[0].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_3 \address_gen[12].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[12].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_2 \address_gen[11].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[11].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_1 \address_gen[10].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[10].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_24 \address_gen[9].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[9].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_23 \address_gen[8].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[8].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_22 \address_gen[7].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[7].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_21 \address_gen[6].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[6].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_20 \address_gen[5].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[5].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_19 \address_gen[4].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[4].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_13 \address_gen[21].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[21].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_12 \address_gen[20].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[20].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_10 \address_gen[19].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[19].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_9 \address_gen[18].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[18].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_8 \address_gen[17].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[17].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_7 \address_gen[16].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[16].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_6 \address_gen[15].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[15].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_5 \address_gen[14].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[14].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_4 \address_gen[13].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[13].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_altddio_out_1 \clock_gen[0].umem_ck_pad (
	.dataout({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }),
	.datain_h({phy_ddio_ck_0}),
	.datain_l({phy_ddio_ck_1}),
	.outclock(\mem_ck_source[0] ));

soc_system_hps_sdram_p0_generic_ddio_3 ureset_n_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk}),
	.dataout({dataout_unconnected_wire_14,dataout_unconnected_wire_13,dataout_unconnected_wire_12,dataout_unconnected_wire_11,dataout_unconnected_wire_10,dataout_unconnected_wire_9,dataout_unconnected_wire_8,dataout_unconnected_wire_7,dataout_unconnected_wire_6,
dataout_unconnected_wire_5,dataout_unconnected_wire_4,dataout_unconnected_wire_3,dataout_unconnected_wire_2,dataout_unconnected_wire_1,dataout_03}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[24].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_reset_n_3,phy_ddio_reset_n_2,phy_ddio_reset_n_1,phy_ddio_reset_n_0}));

soc_system_hps_sdram_p0_generic_ddio_2 ucmd_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_1,dataout_unconnected_wire_13_1,dataout_unconnected_wire_12_1,dataout_unconnected_wire_11_1,dataout_unconnected_wire_10_1,dataout_unconnected_wire_9_1,dataout_unconnected_wire_8_1,dataout_unconnected_wire_7_1,
dataout_unconnected_wire_6_1,dataout_51,dataout_41,dataout_31,dataout_22,dataout_16,dataout_02}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[23].acv_ac_ldc|adc_clk_cps ,\address_gen[22].acv_ac_ldc|adc_clk_cps ,\address_gen[21].acv_ac_ldc|adc_clk_cps ,\address_gen[20].acv_ac_ldc|adc_clk_cps ,\address_gen[19].acv_ac_ldc|adc_clk_cps ,
\address_gen[18].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_we_n_3,phy_ddio_we_n_2,phy_ddio_we_n_1,phy_ddio_we_n_0,phy_ddio_cas_n_3,phy_ddio_cas_n_2,phy_ddio_cas_n_1,phy_ddio_cas_n_0,phy_ddio_ras_n_3,
phy_ddio_ras_n_2,phy_ddio_ras_n_1,phy_ddio_ras_n_0,phy_ddio_odt_3,phy_ddio_odt_2,phy_ddio_odt_1,phy_ddio_odt_0,phy_ddio_cke_3,phy_ddio_cke_2,phy_ddio_cke_1,phy_ddio_cke_0,phy_ddio_cs_n_3,phy_ddio_cs_n_2,phy_ddio_cs_n_1,phy_ddio_cs_n_0}));

soc_system_hps_sdram_p0_generic_ddio_1 ubank_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_2,dataout_unconnected_wire_13_2,dataout_unconnected_wire_12_2,dataout_unconnected_wire_11_2,dataout_unconnected_wire_10_2,dataout_unconnected_wire_9_2,dataout_unconnected_wire_8_2,dataout_unconnected_wire_7_2,
dataout_unconnected_wire_6_2,dataout_unconnected_wire_5_1,dataout_unconnected_wire_4_1,dataout_unconnected_wire_3_1,dataout_21,dataout_15,dataout_01}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[17].acv_ac_ldc|adc_clk_cps ,\address_gen[16].acv_ac_ldc|adc_clk_cps ,\address_gen[15].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_bank_11,phy_ddio_bank_10,phy_ddio_bank_9,phy_ddio_bank_8,phy_ddio_bank_7,phy_ddio_bank_6,phy_ddio_bank_5,
phy_ddio_bank_4,phy_ddio_bank_3,phy_ddio_bank_2,phy_ddio_bank_1,phy_ddio_bank_0}));

soc_system_hps_sdram_p0_generic_ddio uaddress_pad(
	.clk_hr({afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_14,dataout_13,dataout_12,dataout_11,dataout_10,dataout_9,dataout_8,dataout_7,dataout_6,dataout_5,dataout_4,dataout_3,dataout_2,dataout_1,dataout_0}),
	.clk_fr({\address_gen[14].acv_ac_ldc|adc_clk_cps ,\address_gen[13].acv_ac_ldc|adc_clk_cps ,\address_gen[12].acv_ac_ldc|adc_clk_cps ,\address_gen[11].acv_ac_ldc|adc_clk_cps ,\address_gen[10].acv_ac_ldc|adc_clk_cps ,\address_gen[9].acv_ac_ldc|adc_clk_cps ,
\address_gen[8].acv_ac_ldc|adc_clk_cps ,\address_gen[7].acv_ac_ldc|adc_clk_cps ,\address_gen[6].acv_ac_ldc|adc_clk_cps ,\address_gen[5].acv_ac_ldc|adc_clk_cps ,\address_gen[4].acv_ac_ldc|adc_clk_cps ,\address_gen[3].acv_ac_ldc|adc_clk_cps ,
\address_gen[2].acv_ac_ldc|adc_clk_cps ,\address_gen[1].acv_ac_ldc|adc_clk_cps ,\address_gen[0].acv_ac_ldc|adc_clk_cps }),
	.datain({phy_ddio_address_59,phy_ddio_address_58,phy_ddio_address_57,phy_ddio_address_56,phy_ddio_address_55,phy_ddio_address_54,phy_ddio_address_53,phy_ddio_address_52,phy_ddio_address_51,phy_ddio_address_50,phy_ddio_address_49,phy_ddio_address_48,phy_ddio_address_47,
phy_ddio_address_46,phy_ddio_address_45,phy_ddio_address_44,phy_ddio_address_43,phy_ddio_address_42,phy_ddio_address_41,phy_ddio_address_40,phy_ddio_address_39,phy_ddio_address_38,phy_ddio_address_37,phy_ddio_address_36,phy_ddio_address_35,phy_ddio_address_34,
phy_ddio_address_33,phy_ddio_address_32,phy_ddio_address_31,phy_ddio_address_30,phy_ddio_address_29,phy_ddio_address_28,phy_ddio_address_27,phy_ddio_address_26,phy_ddio_address_25,phy_ddio_address_24,phy_ddio_address_23,phy_ddio_address_22,phy_ddio_address_21,
phy_ddio_address_20,phy_ddio_address_19,phy_ddio_address_18,phy_ddio_address_17,phy_ddio_address_16,phy_ddio_address_15,phy_ddio_address_14,phy_ddio_address_13,phy_ddio_address_12,phy_ddio_address_11,phy_ddio_address_10,phy_ddio_address_9,phy_ddio_address_8,
phy_ddio_address_7,phy_ddio_address_6,phy_ddio_address_5,phy_ddio_address_4,phy_ddio_address_3,phy_ddio_address_2,phy_ddio_address_1,phy_ddio_address_0}));

soc_system_hps_sdram_p0_acv_ldc_16 \address_gen[24].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[24].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_15 \address_gen[23].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[23].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_acv_ldc_14 \address_gen[22].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[22].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

soc_system_hps_sdram_p0_clock_pair_generator \clock_gen[0].uclk_generator (
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.datain({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }));

cyclonev_clk_phase_select \clock_gen[0].clk_phase_select_dqs (
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\clock_gen[0].leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(\mem_ck_source[0] ));
defparam \clock_gen[0].clk_phase_select_dqs .invert_phase = "false";
defparam \clock_gen[0].clk_phase_select_dqs .phase_setting = 0;
defparam \clock_gen[0].clk_phase_select_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].clk_phase_select_dqs .use_dqs_input = "false";
defparam \clock_gen[0].clk_phase_select_dqs .use_phasectrlin = "false";

cyclonev_leveling_delay_chain \clock_gen[0].leveling_delay_chain_dqs (
	.clkin(afi_clk),
	.delayctrlin({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.clkout(\clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ));
defparam \clock_gen[0].leveling_delay_chain_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_delay_increment = 10;
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_altddio_out_1 (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
inout 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_ddio_out_uqe auto_generated(
	.dataout({dataout[0]}),
	.datain_h({datain_h[0]}),
	.datain_l({datain_l[0]}),
	.outclock(outclock));

endmodule

module soc_system_ddio_out_uqe (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
output 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "none";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_acv_ldc (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_1 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_2 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_3 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_4 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_5 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_6 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_7 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_8 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_9 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_10 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_11 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_12 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_13 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_14 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_15 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_16 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_17 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_18 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_19 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_20 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_21 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_22 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_23 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_acv_ldc_24 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_p0_clock_pair_generator (
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	datain)/* synthesis synthesis_greybox=0 */;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(datain[0]),
	.oein(gnd),
	.dtcin(gnd),
	.o(wire_pseudo_diffa_o_0),
	.obar(wire_pseudo_diffa_obar_0),
	.oeout(wire_pseudo_diffa_oeout_0),
	.oebout(wire_pseudo_diffa_oebout_0),
	.dtc(),
	.dtcbar());

endmodule

module soc_system_hps_sdram_p0_generic_ddio (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[6].fr_data_lo ;
wire \acblock[6].fr_data_hi ;
wire \acblock[7].fr_data_lo ;
wire \acblock[7].fr_data_hi ;
wire \acblock[8].fr_data_lo ;
wire \acblock[8].fr_data_hi ;
wire \acblock[9].fr_data_lo ;
wire \acblock[9].fr_data_hi ;
wire \acblock[10].fr_data_lo ;
wire \acblock[10].fr_data_hi ;
wire \acblock[11].fr_data_lo ;
wire \acblock[11].fr_data_hi ;
wire \acblock[12].fr_data_lo ;
wire \acblock[12].fr_data_hi ;
wire \acblock[13].fr_data_lo ;
wire \acblock[13].fr_data_hi ;
wire \acblock[14].fr_data_lo ;
wire \acblock[14].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].ddio_out (
	.datainlo(\acblock[6].fr_data_lo ),
	.datainhi(\acblock[6].fr_data_hi ),
	.clkhi(clk_fr[6]),
	.clklo(clk_fr[6]),
	.muxsel(clk_fr[6]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[6]),
	.dfflo(),
	.dffhi());
defparam \acblock[6].ddio_out .async_mode = "none";
defparam \acblock[6].ddio_out .half_rate_mode = "false";
defparam \acblock[6].ddio_out .power_up = "low";
defparam \acblock[6].ddio_out .sync_mode = "none";
defparam \acblock[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].ddio_out (
	.datainlo(\acblock[7].fr_data_lo ),
	.datainhi(\acblock[7].fr_data_hi ),
	.clkhi(clk_fr[7]),
	.clklo(clk_fr[7]),
	.muxsel(clk_fr[7]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[7]),
	.dfflo(),
	.dffhi());
defparam \acblock[7].ddio_out .async_mode = "none";
defparam \acblock[7].ddio_out .half_rate_mode = "false";
defparam \acblock[7].ddio_out .power_up = "low";
defparam \acblock[7].ddio_out .sync_mode = "none";
defparam \acblock[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].ddio_out (
	.datainlo(\acblock[8].fr_data_lo ),
	.datainhi(\acblock[8].fr_data_hi ),
	.clkhi(clk_fr[8]),
	.clklo(clk_fr[8]),
	.muxsel(clk_fr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[8]),
	.dfflo(),
	.dffhi());
defparam \acblock[8].ddio_out .async_mode = "none";
defparam \acblock[8].ddio_out .half_rate_mode = "false";
defparam \acblock[8].ddio_out .power_up = "low";
defparam \acblock[8].ddio_out .sync_mode = "none";
defparam \acblock[8].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].ddio_out (
	.datainlo(\acblock[9].fr_data_lo ),
	.datainhi(\acblock[9].fr_data_hi ),
	.clkhi(clk_fr[9]),
	.clklo(clk_fr[9]),
	.muxsel(clk_fr[9]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[9]),
	.dfflo(),
	.dffhi());
defparam \acblock[9].ddio_out .async_mode = "none";
defparam \acblock[9].ddio_out .half_rate_mode = "false";
defparam \acblock[9].ddio_out .power_up = "low";
defparam \acblock[9].ddio_out .sync_mode = "none";
defparam \acblock[9].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].ddio_out (
	.datainlo(\acblock[10].fr_data_lo ),
	.datainhi(\acblock[10].fr_data_hi ),
	.clkhi(clk_fr[10]),
	.clklo(clk_fr[10]),
	.muxsel(clk_fr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[10]),
	.dfflo(),
	.dffhi());
defparam \acblock[10].ddio_out .async_mode = "none";
defparam \acblock[10].ddio_out .half_rate_mode = "false";
defparam \acblock[10].ddio_out .power_up = "low";
defparam \acblock[10].ddio_out .sync_mode = "none";
defparam \acblock[10].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].ddio_out (
	.datainlo(\acblock[11].fr_data_lo ),
	.datainhi(\acblock[11].fr_data_hi ),
	.clkhi(clk_fr[11]),
	.clklo(clk_fr[11]),
	.muxsel(clk_fr[11]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[11]),
	.dfflo(),
	.dffhi());
defparam \acblock[11].ddio_out .async_mode = "none";
defparam \acblock[11].ddio_out .half_rate_mode = "false";
defparam \acblock[11].ddio_out .power_up = "low";
defparam \acblock[11].ddio_out .sync_mode = "none";
defparam \acblock[11].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].ddio_out (
	.datainlo(\acblock[12].fr_data_lo ),
	.datainhi(\acblock[12].fr_data_hi ),
	.clkhi(clk_fr[12]),
	.clklo(clk_fr[12]),
	.muxsel(clk_fr[12]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[12]),
	.dfflo(),
	.dffhi());
defparam \acblock[12].ddio_out .async_mode = "none";
defparam \acblock[12].ddio_out .half_rate_mode = "false";
defparam \acblock[12].ddio_out .power_up = "low";
defparam \acblock[12].ddio_out .sync_mode = "none";
defparam \acblock[12].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].ddio_out (
	.datainlo(\acblock[13].fr_data_lo ),
	.datainhi(\acblock[13].fr_data_hi ),
	.clkhi(clk_fr[13]),
	.clklo(clk_fr[13]),
	.muxsel(clk_fr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[13]),
	.dfflo(),
	.dffhi());
defparam \acblock[13].ddio_out .async_mode = "none";
defparam \acblock[13].ddio_out .half_rate_mode = "false";
defparam \acblock[13].ddio_out .power_up = "low";
defparam \acblock[13].ddio_out .sync_mode = "none";
defparam \acblock[13].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].ddio_out (
	.datainlo(\acblock[14].fr_data_lo ),
	.datainhi(\acblock[14].fr_data_hi ),
	.clkhi(clk_fr[14]),
	.clklo(clk_fr[14]),
	.muxsel(clk_fr[14]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[14]),
	.dfflo(),
	.dffhi());
defparam \acblock[14].ddio_out .async_mode = "none";
defparam \acblock[14].ddio_out .half_rate_mode = "false";
defparam \acblock[14].ddio_out .power_up = "low";
defparam \acblock[14].ddio_out .sync_mode = "none";
defparam \acblock[14].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_lo (
	.datainlo(datain[27]),
	.datainhi(datain[25]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_lo .async_mode = "none";
defparam \acblock[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_lo .power_up = "low";
defparam \acblock[6].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_hi (
	.datainlo(datain[26]),
	.datainhi(datain[24]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_hi .async_mode = "none";
defparam \acblock[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_hi .power_up = "low";
defparam \acblock[6].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_lo (
	.datainlo(datain[31]),
	.datainhi(datain[29]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_lo .async_mode = "none";
defparam \acblock[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_lo .power_up = "low";
defparam \acblock[7].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_hi (
	.datainlo(datain[30]),
	.datainhi(datain[28]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_hi .async_mode = "none";
defparam \acblock[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_hi .power_up = "low";
defparam \acblock[7].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_lo (
	.datainlo(datain[35]),
	.datainhi(datain[33]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_lo .async_mode = "none";
defparam \acblock[8].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_lo .power_up = "low";
defparam \acblock[8].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[8].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_hi (
	.datainlo(datain[34]),
	.datainhi(datain[32]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_hi .async_mode = "none";
defparam \acblock[8].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_hi .power_up = "low";
defparam \acblock[8].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[8].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_lo (
	.datainlo(datain[39]),
	.datainhi(datain[37]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_lo .async_mode = "none";
defparam \acblock[9].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_lo .power_up = "low";
defparam \acblock[9].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[9].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_hi (
	.datainlo(datain[38]),
	.datainhi(datain[36]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_hi .async_mode = "none";
defparam \acblock[9].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_hi .power_up = "low";
defparam \acblock[9].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[9].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_lo (
	.datainlo(datain[43]),
	.datainhi(datain[41]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_lo .async_mode = "none";
defparam \acblock[10].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_lo .power_up = "low";
defparam \acblock[10].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[10].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_hi (
	.datainlo(datain[42]),
	.datainhi(datain[40]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_hi .async_mode = "none";
defparam \acblock[10].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_hi .power_up = "low";
defparam \acblock[10].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[10].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_lo (
	.datainlo(datain[47]),
	.datainhi(datain[45]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_lo .async_mode = "none";
defparam \acblock[11].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_lo .power_up = "low";
defparam \acblock[11].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[11].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_hi (
	.datainlo(datain[46]),
	.datainhi(datain[44]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_hi .async_mode = "none";
defparam \acblock[11].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_hi .power_up = "low";
defparam \acblock[11].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[11].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_lo (
	.datainlo(datain[51]),
	.datainhi(datain[49]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_lo .async_mode = "none";
defparam \acblock[12].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_lo .power_up = "low";
defparam \acblock[12].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[12].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_hi (
	.datainlo(datain[50]),
	.datainhi(datain[48]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_hi .async_mode = "none";
defparam \acblock[12].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_hi .power_up = "low";
defparam \acblock[12].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[12].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_lo (
	.datainlo(datain[55]),
	.datainhi(datain[53]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_lo .async_mode = "none";
defparam \acblock[13].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_lo .power_up = "low";
defparam \acblock[13].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[13].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_hi (
	.datainlo(datain[54]),
	.datainhi(datain[52]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_hi .async_mode = "none";
defparam \acblock[13].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_hi .power_up = "low";
defparam \acblock[13].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[13].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_lo (
	.datainlo(datain[59]),
	.datainhi(datain[57]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_lo .async_mode = "none";
defparam \acblock[14].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_lo .power_up = "low";
defparam \acblock[14].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[14].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_hi (
	.datainlo(datain[58]),
	.datainhi(datain[56]),
	.clkhi(clk_hr[13]),
	.clklo(clk_hr[13]),
	.muxsel(clk_hr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_hi .async_mode = "none";
defparam \acblock[14].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_hi .power_up = "low";
defparam \acblock[14].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[14].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_generic_ddio_1 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_generic_ddio_2 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[2]),
	.clklo(clk_hr[2]),
	.muxsel(clk_hr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_generic_ddio_3 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_altdqdqs (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_3,phy_ddio_dmdout_2,phy_ddio_dmdout_1,phy_ddio_dmdout_0}),
	.write_data_in({phy_ddio_dqdout_31,phy_ddio_dqdout_30,phy_ddio_dqdout_29,phy_ddio_dqdout_28,phy_ddio_dqdout_27,phy_ddio_dqdout_26,phy_ddio_dqdout_25,phy_ddio_dqdout_24,phy_ddio_dqdout_23,phy_ddio_dqdout_22,phy_ddio_dqdout_21,phy_ddio_dqdout_20,phy_ddio_dqdout_19,phy_ddio_dqdout_18,
phy_ddio_dqdout_17,phy_ddio_dqdout_16,phy_ddio_dqdout_15,phy_ddio_dqdout_14,phy_ddio_dqdout_13,phy_ddio_dqdout_12,phy_ddio_dqdout_11,phy_ddio_dqdout_10,phy_ddio_dqdout_9,phy_ddio_dqdout_8,phy_ddio_dqdout_7,phy_ddio_dqdout_6,phy_ddio_dqdout_5,phy_ddio_dqdout_4,
phy_ddio_dqdout_3,phy_ddio_dqdout_2,phy_ddio_dqdout_1,phy_ddio_dqdout_0}),
	.write_oe_in({phy_ddio_dqoe_15,phy_ddio_dqoe_14,phy_ddio_dqoe_13,phy_ddio_dqoe_12,phy_ddio_dqoe_11,phy_ddio_dqoe_10,phy_ddio_dqoe_9,phy_ddio_dqoe_8,phy_ddio_dqoe_7,phy_ddio_dqoe_6,phy_ddio_dqoe_5,phy_ddio_dqoe_4,phy_ddio_dqoe_3,phy_ddio_dqoe_2,phy_ddio_dqoe_1,phy_ddio_dqoe_0}),
	.write_strobe({phy_ddio_dqs_dout_3,phy_ddio_dqs_dout_2,phy_ddio_dqs_dout_1,phy_ddio_dqs_dout_0}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_0),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_0),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_1,phy_ddio_dqslogic_incrdataen_0}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_1,phy_ddio_dqslogic_incwrptr_0}),
	.oct_ena_in({phy_ddio_dqslogic_oct_1,phy_ddio_dqslogic_oct_0}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_4,phy_ddio_dqslogic_readlatency_3,phy_ddio_dqslogic_readlatency_2,phy_ddio_dqslogic_readlatency_1,phy_ddio_dqslogic_readlatency_0}),
	.output_strobe_ena({phy_ddio_dqs_oe_1,phy_ddio_dqs_oe_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	hr_clock_in,
	write_strobe_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(hr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(hr_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_altdqdqs_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_7,phy_ddio_dmdout_6,phy_ddio_dmdout_5,phy_ddio_dmdout_4}),
	.write_data_in({phy_ddio_dqdout_67,phy_ddio_dqdout_66,phy_ddio_dqdout_65,phy_ddio_dqdout_64,phy_ddio_dqdout_63,phy_ddio_dqdout_62,phy_ddio_dqdout_61,phy_ddio_dqdout_60,phy_ddio_dqdout_59,phy_ddio_dqdout_58,phy_ddio_dqdout_57,phy_ddio_dqdout_56,phy_ddio_dqdout_55,phy_ddio_dqdout_54,
phy_ddio_dqdout_53,phy_ddio_dqdout_52,phy_ddio_dqdout_51,phy_ddio_dqdout_50,phy_ddio_dqdout_49,phy_ddio_dqdout_48,phy_ddio_dqdout_47,phy_ddio_dqdout_46,phy_ddio_dqdout_45,phy_ddio_dqdout_44,phy_ddio_dqdout_43,phy_ddio_dqdout_42,phy_ddio_dqdout_41,phy_ddio_dqdout_40,
phy_ddio_dqdout_39,phy_ddio_dqdout_38,phy_ddio_dqdout_37,phy_ddio_dqdout_36}),
	.write_oe_in({phy_ddio_dqoe_33,phy_ddio_dqoe_32,phy_ddio_dqoe_31,phy_ddio_dqoe_30,phy_ddio_dqoe_29,phy_ddio_dqoe_28,phy_ddio_dqoe_27,phy_ddio_dqoe_26,phy_ddio_dqoe_25,phy_ddio_dqoe_24,phy_ddio_dqoe_23,phy_ddio_dqoe_22,phy_ddio_dqoe_21,phy_ddio_dqoe_20,phy_ddio_dqoe_19,phy_ddio_dqoe_18}),
	.write_strobe({phy_ddio_dqs_dout_7,phy_ddio_dqs_dout_6,phy_ddio_dqs_dout_5,phy_ddio_dqs_dout_4}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_1),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_1),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_3,phy_ddio_dqslogic_incrdataen_2}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_3,phy_ddio_dqslogic_incwrptr_2}),
	.oct_ena_in({phy_ddio_dqslogic_oct_3,phy_ddio_dqslogic_oct_2}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_9,phy_ddio_dqslogic_readlatency_8,phy_ddio_dqslogic_readlatency_7,phy_ddio_dqslogic_readlatency_6,phy_ddio_dqslogic_readlatency_5}),
	.output_strobe_ena({phy_ddio_dqs_oe_3,phy_ddio_dqs_oe_2}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	hr_clock_in,
	write_strobe_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(hr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(hr_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_altdqdqs_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_11,phy_ddio_dmdout_10,phy_ddio_dmdout_9,phy_ddio_dmdout_8}),
	.write_data_in({phy_ddio_dqdout_103,phy_ddio_dqdout_102,phy_ddio_dqdout_101,phy_ddio_dqdout_100,phy_ddio_dqdout_99,phy_ddio_dqdout_98,phy_ddio_dqdout_97,phy_ddio_dqdout_96,phy_ddio_dqdout_95,phy_ddio_dqdout_94,phy_ddio_dqdout_93,phy_ddio_dqdout_92,phy_ddio_dqdout_91,phy_ddio_dqdout_90,
phy_ddio_dqdout_89,phy_ddio_dqdout_88,phy_ddio_dqdout_87,phy_ddio_dqdout_86,phy_ddio_dqdout_85,phy_ddio_dqdout_84,phy_ddio_dqdout_83,phy_ddio_dqdout_82,phy_ddio_dqdout_81,phy_ddio_dqdout_80,phy_ddio_dqdout_79,phy_ddio_dqdout_78,phy_ddio_dqdout_77,phy_ddio_dqdout_76,
phy_ddio_dqdout_75,phy_ddio_dqdout_74,phy_ddio_dqdout_73,phy_ddio_dqdout_72}),
	.write_oe_in({phy_ddio_dqoe_51,phy_ddio_dqoe_50,phy_ddio_dqoe_49,phy_ddio_dqoe_48,phy_ddio_dqoe_47,phy_ddio_dqoe_46,phy_ddio_dqoe_45,phy_ddio_dqoe_44,phy_ddio_dqoe_43,phy_ddio_dqoe_42,phy_ddio_dqoe_41,phy_ddio_dqoe_40,phy_ddio_dqoe_39,phy_ddio_dqoe_38,phy_ddio_dqoe_37,phy_ddio_dqoe_36}),
	.write_strobe({phy_ddio_dqs_dout_11,phy_ddio_dqs_dout_10,phy_ddio_dqs_dout_9,phy_ddio_dqs_dout_8}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_2),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_2),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_5,phy_ddio_dqslogic_incrdataen_4}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_5,phy_ddio_dqslogic_incwrptr_4}),
	.oct_ena_in({phy_ddio_dqslogic_oct_5,phy_ddio_dqslogic_oct_4}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_14,phy_ddio_dqslogic_readlatency_13,phy_ddio_dqslogic_readlatency_12,phy_ddio_dqslogic_readlatency_11,phy_ddio_dqslogic_readlatency_10}),
	.output_strobe_ena({phy_ddio_dqs_oe_5,phy_ddio_dqs_oe_4}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	hr_clock_in,
	write_strobe_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(hr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(hr_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_altdqdqs_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.config_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_15,phy_ddio_dmdout_14,phy_ddio_dmdout_13,phy_ddio_dmdout_12}),
	.write_data_in({phy_ddio_dqdout_139,phy_ddio_dqdout_138,phy_ddio_dqdout_137,phy_ddio_dqdout_136,phy_ddio_dqdout_135,phy_ddio_dqdout_134,phy_ddio_dqdout_133,phy_ddio_dqdout_132,phy_ddio_dqdout_131,phy_ddio_dqdout_130,phy_ddio_dqdout_129,phy_ddio_dqdout_128,phy_ddio_dqdout_127,
phy_ddio_dqdout_126,phy_ddio_dqdout_125,phy_ddio_dqdout_124,phy_ddio_dqdout_123,phy_ddio_dqdout_122,phy_ddio_dqdout_121,phy_ddio_dqdout_120,phy_ddio_dqdout_119,phy_ddio_dqdout_118,phy_ddio_dqdout_117,phy_ddio_dqdout_116,phy_ddio_dqdout_115,phy_ddio_dqdout_114,
phy_ddio_dqdout_113,phy_ddio_dqdout_112,phy_ddio_dqdout_111,phy_ddio_dqdout_110,phy_ddio_dqdout_109,phy_ddio_dqdout_108}),
	.write_oe_in({phy_ddio_dqoe_69,phy_ddio_dqoe_68,phy_ddio_dqoe_67,phy_ddio_dqoe_66,phy_ddio_dqoe_65,phy_ddio_dqoe_64,phy_ddio_dqoe_63,phy_ddio_dqoe_62,phy_ddio_dqoe_61,phy_ddio_dqoe_60,phy_ddio_dqoe_59,phy_ddio_dqoe_58,phy_ddio_dqoe_57,phy_ddio_dqoe_56,phy_ddio_dqoe_55,phy_ddio_dqoe_54}),
	.write_strobe({phy_ddio_dqs_dout_15,phy_ddio_dqs_dout_14,phy_ddio_dqs_dout_13,phy_ddio_dqs_dout_12}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_3),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_3),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_7,phy_ddio_dqslogic_incrdataen_6}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_7,phy_ddio_dqslogic_incwrptr_6}),
	.oct_ena_in({phy_ddio_dqslogic_oct_7,phy_ddio_dqslogic_oct_6}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_19,phy_ddio_dqslogic_readlatency_18,phy_ddio_dqslogic_readlatency_17,phy_ddio_dqslogic_readlatency_16,phy_ddio_dqslogic_readlatency_15}),
	.output_strobe_ena({phy_ddio_dqs_oe_7,phy_ddio_dqs_oe_6}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module soc_system_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	hr_clock_in,
	write_strobe_clock_in,
	config_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	vfifo_qvld,
	lfifo_rdata_en_full,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	config_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] vfifo_qvld;
input 	[1:0] lfifo_rdata_en_full;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(hr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(hr_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(hr_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(vfifo_qvld[1]),
	.datainhi(vfifo_qvld[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module soc_system_hps_sdram_p0_acv_ldc_25 (
	pll_hr_clk,
	pll_dqs_clk,
	adc_clk,
	avl_clk,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_hr_clk;
input 	pll_dqs_clk;
output 	adc_clk;
output 	avl_clk;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;

assign adc_clk = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

assign avl_clk = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_hr_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(pll_hr_clk),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

endmodule

module soc_system_hps_sdram_pll (
	afi_half_clk,
	pll_write_clk_pre_phy_clk)/* synthesis synthesis_greybox=0 */;
output 	afi_half_clk;
output 	pll_write_clk_pre_phy_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_out[2] ;
wire \clk_out[3] ;

wire [3:0] pll_CLK_OUT_bus;

assign afi_half_clk = pll_CLK_OUT_bus[0];
assign pll_write_clk_pre_phy_clk = pll_CLK_OUT_bus[1];
assign \clk_out[2]  = pll_CLK_OUT_bus[2];
assign \clk_out[3]  = pll_CLK_OUT_bus[3];

cyclonev_hps_sdram_pll pll(
	.ref_clk(gnd),
	.clk_out(pll_CLK_OUT_bus));

endmodule

module soc_system_soc_system_mm_interconnect_0 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	source0_data_34,
	source0_data_32,
	sink1_ready,
	hps_0_h2f_lw_axi_master_awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	hps_0_h2f_lw_axi_master_wready,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	int_nxt_addr_reg_dly_10,
	int_nxt_addr_reg_dly_11,
	int_nxt_addr_reg_dly_12,
	int_nxt_addr_reg_dly_13,
	int_nxt_addr_reg_dly_14,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	source0_data_33,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	source0_data_35,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	altera_reset_synchronizer_int_chain_out,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARADDR_6;
input 	h2f_lw_ARADDR_7;
input 	h2f_lw_ARADDR_8;
input 	h2f_lw_ARADDR_9;
input 	h2f_lw_ARADDR_10;
input 	h2f_lw_ARADDR_11;
input 	h2f_lw_ARADDR_12;
input 	h2f_lw_ARADDR_13;
input 	h2f_lw_ARADDR_14;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_17;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
output 	source0_data_34;
output 	source0_data_32;
output 	sink1_ready;
output 	hps_0_h2f_lw_axi_master_awready;
output 	src0_valid;
output 	source_endofpacket;
output 	src1_valid;
output 	hps_0_h2f_lw_axi_master_wready;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	out_data_19;
output 	out_data_20;
output 	out_data_21;
output 	out_data_22;
output 	out_data_23;
output 	out_data_24;
output 	out_data_25;
output 	out_data_26;
output 	out_data_27;
output 	out_data_28;
output 	out_data_29;
output 	out_data_30;
output 	out_data_31;
output 	m0_write;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
output 	int_nxt_addr_reg_dly_10;
output 	int_nxt_addr_reg_dly_11;
output 	int_nxt_addr_reg_dly_12;
output 	int_nxt_addr_reg_dly_13;
output 	int_nxt_addr_reg_dly_14;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	source0_data_33;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	source0_data_35;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	altera_reset_synchronizer_int_chain_out;
input 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~21_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~21_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ;
wire \hps_0_h2f_lw_axi_master_agent|Add5~25_sumout ;
wire \hps_0_h2f_lw_axi_master_agent|Add4~25_sumout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~6_combout ;
wire \onchip_memory2_0_s1_agent|WideOr0~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ;
wire \cmd_mux|saved_grant[0]~q ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_memory2_0_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][112]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \onchip_memory2_0_s1_agent|uncompressor|always0~0_combout ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][59]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux|src0_valid~0_combout ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][113]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \onchip_memory2_0_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \cmd_mux|src_valid~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \onchip_memory2_0_s1_agent|m0_write~0_combout ;
wire \cmd_mux|WideOr1~combout ;
wire \cmd_mux|src_payload[0]~combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \hps_0_h2f_lw_axi_master_agent|sop_enable~q ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[6]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ;
wire \hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ;
wire \hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~4_combout ;
wire \onchip_memory2_0_s1_agent|comb~0_combout ;
wire \rsp_demux|WideOr0~0_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \cmd_mux|src_data[78]~combout ;
wire \cmd_mux|src_data[79]~combout ;
wire \cmd_mux|src_data[77]~combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add1~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|log2ceil~0_combout ;
wire \cmd_mux|src_payload~2_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add3~0_combout ;
wire \hps_0_h2f_lw_axi_master_agent|log2ceil~1_combout ;
wire \cmd_mux|src_data[71]~3_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~0_combout ;
wire \cmd_mux|src_payload~4_combout ;
wire \hps_0_h2f_lw_axi_master_agent|log2ceil~2_combout ;
wire \cmd_mux|src_payload~5_combout ;
wire \hps_0_h2f_lw_axi_master_agent|Add3~1_combout ;
wire \cmd_mux|src_data[70]~6_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~1_combout ;
wire \cmd_mux|src_data[34]~combout ;
wire \cmd_mux|src_data[32]~combout ;
wire \cmd_mux|src_data[35]~combout ;
wire \cmd_mux|src_data[33]~combout ;
wire \onchip_memory2_0_s1_agent|cp_ready~1_combout ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \cmd_mux|src_payload~6_combout ;
wire \cmd_mux|src_payload~7_combout ;
wire \cmd_mux|src_payload~8_combout ;
wire \cmd_mux|src_data[72]~9_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~2_combout ;
wire \cmd_mux|src_payload~9_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ;
wire \cmd_mux|src_data[73]~11_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~3_combout ;
wire \cmd_mux|src_payload~10_combout ;
wire \cmd_mux|src_payload~11_combout ;
wire \cmd_mux|src_data[74]~13_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~4_combout ;
wire \cmd_mux|src_payload~12_combout ;
wire \cmd_mux|src_payload~13_combout ;
wire \cmd_mux|src_data[75]~15_combout ;
wire \hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~5_combout ;
wire \cmd_mux|src_payload~14_combout ;
wire \cmd_mux|src_payload~15_combout ;
wire \cmd_mux|src_payload~16_combout ;
wire \cmd_mux|src_payload~17_combout ;
wire \cmd_mux|src_payload~18_combout ;
wire \cmd_mux|src_payload~19_combout ;
wire \cmd_mux|src_payload~20_combout ;
wire \cmd_mux|src_payload~21_combout ;
wire \cmd_mux|src_payload~22_combout ;
wire \cmd_mux|src_payload~23_combout ;
wire \cmd_mux|src_payload~24_combout ;
wire \cmd_mux|src_payload~25_combout ;
wire \cmd_mux|src_payload~26_combout ;
wire \cmd_mux|src_payload~27_combout ;
wire \cmd_mux|src_payload~28_combout ;
wire \cmd_mux|src_payload~29_combout ;
wire \cmd_mux|src_payload~30_combout ;
wire \cmd_mux|src_payload~31_combout ;
wire \cmd_mux|src_payload~32_combout ;
wire \cmd_mux|src_payload~33_combout ;
wire \cmd_mux|src_payload~34_combout ;
wire \cmd_mux|src_payload~35_combout ;
wire \cmd_mux|src_payload~36_combout ;
wire \cmd_mux|src_payload~37_combout ;
wire \cmd_mux|src_payload~38_combout ;
wire \cmd_mux|src_payload~39_combout ;
wire \cmd_mux|src_payload~40_combout ;
wire \cmd_mux|src_payload~41_combout ;
wire \cmd_mux|src_payload~42_combout ;
wire \cmd_mux|src_payload~43_combout ;
wire \cmd_mux|src_payload~44_combout ;
wire \cmd_mux|src_data[71]~16_combout ;
wire \cmd_mux|src_data[70]~17_combout ;
wire \cmd_mux|src_data[88]~combout ;
wire \cmd_mux|src_data[89]~combout ;
wire \cmd_mux|src_data[90]~combout ;
wire \cmd_mux|src_data[91]~combout ;
wire \cmd_mux|src_data[92]~combout ;
wire \cmd_mux|src_data[93]~combout ;
wire \cmd_mux|src_data[94]~combout ;
wire \cmd_mux|src_data[95]~combout ;
wire \cmd_mux|src_data[96]~combout ;
wire \cmd_mux|src_data[97]~combout ;
wire \cmd_mux|src_data[98]~combout ;
wire \cmd_mux|src_data[99]~combout ;
wire \cmd_mux|src_data[72]~18_combout ;
wire \cmd_mux|src_data[73]~19_combout ;
wire \cmd_mux|src_data[74]~20_combout ;
wire \cmd_mux|src_data[75]~21_combout ;
wire \cmd_mux|src_data[76]~22_combout ;
wire \cmd_mux|src_data[76]~23_combout ;
wire \cmd_mux|src_data[76]~25_combout ;


soc_system_soc_system_mm_interconnect_0_rsp_demux rsp_demux(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_memory2_0_s1_agent_rdata_fifo|mem_used[0]~q ),
	.always0(\onchip_memory2_0_s1_agent|uncompressor|always0~0_combout ),
	.mem_59_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux|src0_valid~0_combout ),
	.src0_valid2(src0_valid),
	.src1_valid(src1_valid),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

soc_system_soc_system_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.outclk_wire_0(outclk_wire_0),
	.Add4(\hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add5(\hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add41(\hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add51(\hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add42(\hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add52(\hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add43(\hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add53(\hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add44(\hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.Add54(\hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.Add45(\hps_0_h2f_lw_axi_master_agent|Add4~21_sumout ),
	.Add55(\hps_0_h2f_lw_axi_master_agent|Add5~21_sumout ),
	.Add56(\hps_0_h2f_lw_axi_master_agent|Add5~25_sumout ),
	.Add46(\hps_0_h2f_lw_axi_master_agent|Add4~25_sumout ),
	.nxt_out_eop(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.new_burst_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ),
	.nxt_in_ready(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.sink1_ready1(sink1_ready),
	.nxt_in_ready3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.WideOr11(\cmd_mux|WideOr1~combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.Add1(\hps_0_h2f_lw_axi_master_agent|Add1~0_combout ),
	.log2ceil(\hps_0_h2f_lw_axi_master_agent|log2ceil~0_combout ),
	.src_payload1(\cmd_mux|src_payload~2_combout ),
	.Add3(\hps_0_h2f_lw_axi_master_agent|Add3~0_combout ),
	.log2ceil1(\hps_0_h2f_lw_axi_master_agent|log2ceil~1_combout ),
	.src_data_71(\cmd_mux|src_data[71]~3_combout ),
	.src_payload2(\cmd_mux|src_payload~4_combout ),
	.log2ceil2(\hps_0_h2f_lw_axi_master_agent|log2ceil~2_combout ),
	.src_payload3(\cmd_mux|src_payload~5_combout ),
	.Add31(\hps_0_h2f_lw_axi_master_agent|Add3~1_combout ),
	.src_data_70(\cmd_mux|src_data[70]~6_combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_payload4(\cmd_mux|src_payload~6_combout ),
	.src_payload5(\cmd_mux|src_payload~7_combout ),
	.src_payload6(\cmd_mux|src_payload~8_combout ),
	.src_data_72(\cmd_mux|src_data[72]~9_combout ),
	.src_payload7(\cmd_mux|src_payload~9_combout ),
	.Selector17(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ),
	.src_data_73(\cmd_mux|src_data[73]~11_combout ),
	.src_payload8(\cmd_mux|src_payload~10_combout ),
	.src_payload9(\cmd_mux|src_payload~11_combout ),
	.src_data_74(\cmd_mux|src_data[74]~13_combout ),
	.src_payload10(\cmd_mux|src_payload~12_combout ),
	.src_payload11(\cmd_mux|src_payload~13_combout ),
	.src_data_75(\cmd_mux|src_data[75]~15_combout ),
	.src_payload12(\cmd_mux|src_payload~14_combout ),
	.src_payload13(\cmd_mux|src_payload~15_combout ),
	.src_payload14(\cmd_mux|src_payload~16_combout ),
	.src_payload15(\cmd_mux|src_payload~17_combout ),
	.src_payload16(\cmd_mux|src_payload~18_combout ),
	.src_payload17(\cmd_mux|src_payload~19_combout ),
	.src_payload18(\cmd_mux|src_payload~20_combout ),
	.src_payload19(\cmd_mux|src_payload~21_combout ),
	.src_payload20(\cmd_mux|src_payload~22_combout ),
	.src_payload21(\cmd_mux|src_payload~23_combout ),
	.src_payload22(\cmd_mux|src_payload~24_combout ),
	.src_payload23(\cmd_mux|src_payload~25_combout ),
	.src_payload24(\cmd_mux|src_payload~26_combout ),
	.src_payload25(\cmd_mux|src_payload~27_combout ),
	.src_payload26(\cmd_mux|src_payload~28_combout ),
	.src_payload27(\cmd_mux|src_payload~29_combout ),
	.src_payload28(\cmd_mux|src_payload~30_combout ),
	.src_payload29(\cmd_mux|src_payload~31_combout ),
	.src_payload30(\cmd_mux|src_payload~32_combout ),
	.src_payload31(\cmd_mux|src_payload~33_combout ),
	.src_payload32(\cmd_mux|src_payload~34_combout ),
	.src_payload33(\cmd_mux|src_payload~35_combout ),
	.src_payload34(\cmd_mux|src_payload~36_combout ),
	.src_payload35(\cmd_mux|src_payload~37_combout ),
	.src_payload36(\cmd_mux|src_payload~38_combout ),
	.src_payload37(\cmd_mux|src_payload~39_combout ),
	.src_payload38(\cmd_mux|src_payload~40_combout ),
	.src_payload39(\cmd_mux|src_payload~41_combout ),
	.src_payload40(\cmd_mux|src_payload~42_combout ),
	.src_payload41(\cmd_mux|src_payload~43_combout ),
	.src_payload42(\cmd_mux|src_payload~44_combout ),
	.src_data_711(\cmd_mux|src_data[71]~16_combout ),
	.src_data_701(\cmd_mux|src_data[70]~17_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_data_721(\cmd_mux|src_data[72]~18_combout ),
	.src_data_731(\cmd_mux|src_data[73]~19_combout ),
	.src_data_741(\cmd_mux|src_data[74]~20_combout ),
	.src_data_751(\cmd_mux|src_data[75]~21_combout ),
	.src_data_76(\cmd_mux|src_data[76]~22_combout ),
	.src_data_761(\cmd_mux|src_data[76]~23_combout ),
	.src_data_762(\cmd_mux|src_data[76]~25_combout ));

soc_system_altera_merlin_burst_adapter onchip_memory2_0_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARADDR_5(h2f_lw_ARADDR_5),
	.h2f_lw_ARADDR_6(h2f_lw_ARADDR_6),
	.h2f_lw_ARADDR_7(h2f_lw_ARADDR_7),
	.h2f_lw_ARADDR_8(h2f_lw_ARADDR_8),
	.h2f_lw_ARADDR_9(h2f_lw_ARADDR_9),
	.h2f_lw_ARADDR_10(h2f_lw_ARADDR_10),
	.h2f_lw_ARADDR_11(h2f_lw_ARADDR_11),
	.h2f_lw_ARADDR_12(h2f_lw_ARADDR_12),
	.h2f_lw_ARADDR_13(h2f_lw_ARADDR_13),
	.h2f_lw_ARADDR_14(h2f_lw_ARADDR_14),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.outclk_wire_0(outclk_wire_0),
	.address_burst_6(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_7(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_8(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_9(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_10(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_11(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_12(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.address_burst_13(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_14(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.nxt_out_eop(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.new_burst_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ),
	.mem_used_1(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_ready_hold(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_narrow_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.source0_data_33(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~0_combout ),
	.in_byteen_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.source0_data_32(source0_data_32),
	.source0_data_35(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ),
	.in_byteen_reg_3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.source0_data_351(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ),
	.in_byteen_reg_1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.source0_data_331(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~6_combout ),
	.WideOr0(\onchip_memory2_0_s1_agent|WideOr0~0_combout ),
	.nxt_in_ready(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.nxt_in_ready3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.in_data_reg_59(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_5(int_nxt_addr_reg_dly_5),
	.int_nxt_addr_reg_dly_6(int_nxt_addr_reg_dly_6),
	.int_nxt_addr_reg_dly_7(int_nxt_addr_reg_dly_7),
	.int_nxt_addr_reg_dly_8(int_nxt_addr_reg_dly_8),
	.int_nxt_addr_reg_dly_9(int_nxt_addr_reg_dly_9),
	.int_nxt_addr_reg_dly_10(int_nxt_addr_reg_dly_10),
	.int_nxt_addr_reg_dly_11(int_nxt_addr_reg_dly_11),
	.int_nxt_addr_reg_dly_12(int_nxt_addr_reg_dly_12),
	.int_nxt_addr_reg_dly_13(int_nxt_addr_reg_dly_13),
	.int_nxt_addr_reg_dly_14(int_nxt_addr_reg_dly_14),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.source0_data_332(source0_data_33),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.source0_data_352(source0_data_35),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.WideOr1(\cmd_mux|WideOr1~combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.nxt_out_eop1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.sop_enable(\hps_0_h2f_lw_axi_master_agent|sop_enable~q ),
	.burst_bytecount_6(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.burst_bytecount_5(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_4(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\hps_0_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ),
	.burst_bytecount_3(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~4_combout ),
	.in_data_reg_60(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_data_71(\cmd_mux|src_data[71]~3_combout ),
	.out_data_1(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~0_combout ),
	.src_payload1(\cmd_mux|src_payload~4_combout ),
	.src_data_70(\cmd_mux|src_data[70]~6_combout ),
	.out_data_0(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~1_combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.cp_ready(\onchip_memory2_0_s1_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_5(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_88(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.src_payload2(\cmd_mux|src_payload~6_combout ),
	.src_payload3(\cmd_mux|src_payload~7_combout ),
	.src_data_72(\cmd_mux|src_data[72]~9_combout ),
	.out_data_2(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~2_combout ),
	.src_payload4(\cmd_mux|src_payload~9_combout ),
	.src_data_73(\cmd_mux|src_data[73]~11_combout ),
	.out_data_3(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~3_combout ),
	.src_payload5(\cmd_mux|src_payload~10_combout ),
	.src_data_74(\cmd_mux|src_data[74]~13_combout ),
	.out_data_4(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~4_combout ),
	.src_payload6(\cmd_mux|src_payload~12_combout ),
	.src_data_75(\cmd_mux|src_data[75]~15_combout ),
	.out_data_5(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~5_combout ),
	.src_payload7(\cmd_mux|src_payload~14_combout ),
	.src_payload8(\cmd_mux|src_payload~15_combout ),
	.src_payload9(\cmd_mux|src_payload~16_combout ),
	.src_payload10(\cmd_mux|src_payload~17_combout ),
	.src_payload11(\cmd_mux|src_payload~18_combout ),
	.src_payload12(\cmd_mux|src_payload~19_combout ),
	.src_payload13(\cmd_mux|src_payload~20_combout ),
	.src_payload14(\cmd_mux|src_payload~21_combout ),
	.src_payload15(\cmd_mux|src_payload~22_combout ),
	.src_payload16(\cmd_mux|src_payload~23_combout ),
	.src_payload17(\cmd_mux|src_payload~24_combout ),
	.src_payload18(\cmd_mux|src_payload~25_combout ),
	.src_payload19(\cmd_mux|src_payload~26_combout ),
	.src_payload20(\cmd_mux|src_payload~27_combout ),
	.src_payload21(\cmd_mux|src_payload~28_combout ),
	.src_payload22(\cmd_mux|src_payload~29_combout ),
	.src_payload23(\cmd_mux|src_payload~30_combout ),
	.src_payload24(\cmd_mux|src_payload~31_combout ),
	.src_payload25(\cmd_mux|src_payload~32_combout ),
	.src_payload26(\cmd_mux|src_payload~33_combout ),
	.src_payload27(\cmd_mux|src_payload~34_combout ),
	.src_payload28(\cmd_mux|src_payload~35_combout ),
	.src_payload29(\cmd_mux|src_payload~36_combout ),
	.src_payload30(\cmd_mux|src_payload~37_combout ),
	.src_payload31(\cmd_mux|src_payload~38_combout ),
	.src_payload32(\cmd_mux|src_payload~39_combout ),
	.src_payload33(\cmd_mux|src_payload~40_combout ),
	.src_payload34(\cmd_mux|src_payload~41_combout ),
	.src_payload35(\cmd_mux|src_payload~42_combout ),
	.src_payload36(\cmd_mux|src_payload~43_combout ),
	.src_payload37(\cmd_mux|src_payload~44_combout ),
	.src_data_711(\cmd_mux|src_data[71]~16_combout ),
	.src_data_701(\cmd_mux|src_data[70]~17_combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.src_data_721(\cmd_mux|src_data[72]~18_combout ),
	.src_data_731(\cmd_mux|src_data[73]~19_combout ),
	.src_data_741(\cmd_mux|src_data[74]~20_combout ),
	.src_data_751(\cmd_mux|src_data[75]~21_combout ),
	.src_data_76(\cmd_mux|src_data[76]~22_combout ),
	.src_data_761(\cmd_mux|src_data[76]~23_combout ),
	.src_data_762(\cmd_mux|src_data[76]~25_combout ));

soc_system_altera_avalon_sc_fifo onchip_memory2_0_s1_agent_rdata_fifo(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.clk(outclk_wire_0),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_10(q_a_10),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_16(q_a_16),
	.q_a_17(q_a_17),
	.q_a_18(q_a_18),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.q_a_21(q_a_21),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_memory2_0_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[0]~q ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.out_data_0(out_data_0),
	.out_data_1(out_data_1),
	.out_data_2(out_data_2),
	.out_data_3(out_data_3),
	.out_data_4(out_data_4),
	.out_data_5(out_data_5),
	.out_data_6(out_data_6),
	.out_data_7(out_data_7),
	.out_data_8(out_data_8),
	.out_data_9(out_data_9),
	.out_data_10(out_data_10),
	.out_data_11(out_data_11),
	.out_data_12(out_data_12),
	.out_data_13(out_data_13),
	.out_data_14(out_data_14),
	.out_data_15(out_data_15),
	.out_data_16(out_data_16),
	.out_data_17(out_data_17),
	.out_data_18(out_data_18),
	.out_data_19(out_data_19),
	.out_data_20(out_data_20),
	.out_data_21(out_data_21),
	.out_data_22(out_data_22),
	.out_data_23(out_data_23),
	.out_data_24(out_data_24),
	.out_data_25(out_data_25),
	.out_data_26(out_data_26),
	.out_data_27(out_data_27),
	.out_data_28(out_data_28),
	.out_data_29(out_data_29),
	.out_data_30(out_data_30),
	.out_data_31(out_data_31),
	.reset(altera_reset_synchronizer_int_chain_out));

soc_system_altera_avalon_sc_fifo_1 onchip_memory2_0_s1_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.nxt_out_eop(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.mem_used_1(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_ready_hold(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.source0_data_34(source0_data_34),
	.WideOr0(\onchip_memory2_0_s1_agent|WideOr0~0_combout ),
	.out_valid_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_112_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_113_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_69_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\onchip_memory2_0_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.mem_88_0(mem_88_0),
	.mem_89_0(mem_89_0),
	.mem_90_0(mem_90_0),
	.mem_91_0(mem_91_0),
	.mem_92_0(mem_92_0),
	.mem_93_0(mem_93_0),
	.mem_94_0(mem_94_0),
	.mem_95_0(mem_95_0),
	.mem_96_0(mem_96_0),
	.mem_97_0(mem_97_0),
	.mem_98_0(mem_98_0),
	.mem_99_0(mem_99_0),
	.in_data_reg_59(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.m0_write(\onchip_memory2_0_s1_agent|m0_write~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_byte_cnt_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.comb(\onchip_memory2_0_s1_agent|comb~0_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.in_data_reg_60(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.out_uncomp_byte_cnt_reg_5(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_88(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ));

soc_system_altera_merlin_slave_agent onchip_memory2_0_s1_agent(
	.outclk_wire_0(outclk_wire_0),
	.mem_used_1(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_ready_hold(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_narrow_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.source0_data_33(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~0_combout ),
	.in_byteen_reg_2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.source0_data_32(source0_data_32),
	.source0_data_35(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ),
	.in_byteen_reg_3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.source0_data_351(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ),
	.in_byteen_reg_1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.source0_data_331(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~6_combout ),
	.WideOr0(\onchip_memory2_0_s1_agent|WideOr0~0_combout ),
	.out_valid_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_memory2_0_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\onchip_memory2_0_s1_agent_rsp_fifo|mem_used[0]~q ),
	.always0(\onchip_memory2_0_s1_agent|uncompressor|always0~0_combout ),
	.mem_57_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_113_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][113]~q ),
	.mem_69_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\onchip_memory2_0_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.source_endofpacket(source_endofpacket),
	.in_data_reg_59(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.m0_write(\onchip_memory2_0_s1_agent|m0_write~0_combout ),
	.m0_write1(m0_write),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.comb(\onchip_memory2_0_s1_agent|comb~0_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.cp_ready(\onchip_memory2_0_s1_agent|cp_ready~1_combout ));

soc_system_altera_merlin_axi_master_ni hps_0_h2f_lw_axi_master_agent(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.outclk_wire_0(outclk_wire_0),
	.Add4(\hps_0_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add5(\hps_0_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add41(\hps_0_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add51(\hps_0_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add42(\hps_0_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add52(\hps_0_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add43(\hps_0_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add53(\hps_0_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add44(\hps_0_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.Add54(\hps_0_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.Add45(\hps_0_h2f_lw_axi_master_agent|Add4~21_sumout ),
	.Add55(\hps_0_h2f_lw_axi_master_agent|Add5~21_sumout ),
	.address_burst_6(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_7(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_8(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_9(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_10(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_11(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_12(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.address_burst_13(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_14(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.Add56(\hps_0_h2f_lw_axi_master_agent|Add5~25_sumout ),
	.Add46(\hps_0_h2f_lw_axi_master_agent|Add4~25_sumout ),
	.nxt_out_eop(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.new_burst_reg(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ),
	.nxt_in_ready(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~3_combout ),
	.nxt_in_ready3(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.awready(hps_0_h2f_lw_axi_master_awready),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.wready(hps_0_h2f_lw_axi_master_wready),
	.sop_enable1(\hps_0_h2f_lw_axi_master_agent|sop_enable~q ),
	.burst_bytecount_6(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\hps_0_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.burst_bytecount_5(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\hps_0_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_4(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\hps_0_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_2(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\hps_0_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ),
	.burst_bytecount_3(\hps_0_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\hps_0_h2f_lw_axi_master_agent|write_cp_data[66]~4_combout ),
	.Add1(\hps_0_h2f_lw_axi_master_agent|Add1~0_combout ),
	.log2ceil(\hps_0_h2f_lw_axi_master_agent|log2ceil~0_combout ),
	.src_payload(\cmd_mux|src_payload~2_combout ),
	.Add3(\hps_0_h2f_lw_axi_master_agent|Add3~0_combout ),
	.log2ceil1(\hps_0_h2f_lw_axi_master_agent|log2ceil~1_combout ),
	.out_data_1(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~0_combout ),
	.log2ceil2(\hps_0_h2f_lw_axi_master_agent|log2ceil~2_combout ),
	.src_payload1(\cmd_mux|src_payload~5_combout ),
	.Add31(\hps_0_h2f_lw_axi_master_agent|Add3~1_combout ),
	.out_data_0(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~1_combout ),
	.src_payload2(\cmd_mux|src_payload~8_combout ),
	.out_data_2(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~2_combout ),
	.Selector17(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ),
	.out_data_3(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~3_combout ),
	.src_payload3(\cmd_mux|src_payload~11_combout ),
	.out_data_4(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~4_combout ),
	.src_payload4(\cmd_mux|src_payload~13_combout ),
	.out_data_5(\hps_0_h2f_lw_axi_master_agent|align_address_to_size|out_data[5]~5_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1));

soc_system_altera_merlin_slave_translator onchip_memory2_0_s1_translator(
	.clk(outclk_wire_0),
	.in_ready_hold(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.source0_data_34(source0_data_34),
	.WideOr0(\onchip_memory2_0_s1_agent|WideOr0~0_combout ),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write(\onchip_memory2_0_s1_agent|m0_write~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_60(\onchip_memory2_0_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ));

endmodule

module soc_system_altera_avalon_sc_fifo (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	clk,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	src0_valid,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	reset)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	clk;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_17;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	src0_valid;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	out_data_19;
output 	out_data_20;
output 	out_data_21;
output 	out_data_22;
output 	out_data_23;
output 	out_data_24;
output 	out_data_25;
output 	out_data_26;
output 	out_data_27;
output 	out_data_28;
output 	out_data_29;
output 	out_data_30;
output 	out_data_31;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \read~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[0][2]~q ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[0][3]~q ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[0][4]~q ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[0][5]~q ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[0][6]~q ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[0][7]~q ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[0][8]~q ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[0][9]~q ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[0][10]~q ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[0][11]~q ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[0][12]~q ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[0][13]~q ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[0][14]~q ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[0][15]~q ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[0][16]~q ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[0][17]~q ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[0][18]~q ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[0][19]~q ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[0][20]~q ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[0][21]~q ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[0][22]~q ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[0][23]~q ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[0][24]~q ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[0][25]~q ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[0][26]~q ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[0][27]~q ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[0][28]~q ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[0][29]~q ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[0][30]~q ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;
wire \mem[0][31]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \out_data[0]~0 (
	.dataa(!q_a_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~0 .extended_lut = "off";
defparam \out_data[0]~0 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~1 (
	.dataa(!q_a_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~1 .extended_lut = "off";
defparam \out_data[1]~1 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~2 (
	.dataa(!q_a_2),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~2 .extended_lut = "off";
defparam \out_data[2]~2 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~3 (
	.dataa(!q_a_3),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~3 .extended_lut = "off";
defparam \out_data[3]~3 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~4 (
	.dataa(!q_a_4),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~4 .extended_lut = "off";
defparam \out_data[4]~4 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~5 (
	.dataa(!q_a_5),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~5 .extended_lut = "off";
defparam \out_data[5]~5 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~6 (
	.dataa(!q_a_6),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~6 .extended_lut = "off";
defparam \out_data[6]~6 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~7 (
	.dataa(!q_a_7),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~7 .extended_lut = "off";
defparam \out_data[7]~7 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~8 (
	.dataa(!q_a_8),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~8 .extended_lut = "off";
defparam \out_data[8]~8 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~9 (
	.dataa(!q_a_9),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~9 .extended_lut = "off";
defparam \out_data[9]~9 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[9]~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~10 (
	.dataa(!q_a_10),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~10 .extended_lut = "off";
defparam \out_data[10]~10 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~11 (
	.dataa(!q_a_11),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~11 .extended_lut = "off";
defparam \out_data[11]~11 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~12 (
	.dataa(!q_a_12),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~12 .extended_lut = "off";
defparam \out_data[12]~12 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~13 (
	.dataa(!q_a_13),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~13 .extended_lut = "off";
defparam \out_data[13]~13 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~14 (
	.dataa(!q_a_14),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~14 .extended_lut = "off";
defparam \out_data[14]~14 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[14]~14 .shared_arith = "off";

cyclonev_lcell_comb \out_data[15]~15 (
	.dataa(!q_a_15),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[15]~15 .extended_lut = "off";
defparam \out_data[15]~15 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[15]~15 .shared_arith = "off";

cyclonev_lcell_comb \out_data[16]~16 (
	.dataa(!q_a_16),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[16]~16 .extended_lut = "off";
defparam \out_data[16]~16 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[16]~16 .shared_arith = "off";

cyclonev_lcell_comb \out_data[17]~17 (
	.dataa(!q_a_17),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[17]~17 .extended_lut = "off";
defparam \out_data[17]~17 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[17]~17 .shared_arith = "off";

cyclonev_lcell_comb \out_data[18]~18 (
	.dataa(!q_a_18),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[18]~18 .extended_lut = "off";
defparam \out_data[18]~18 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[18]~18 .shared_arith = "off";

cyclonev_lcell_comb \out_data[19]~19 (
	.dataa(!q_a_19),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[19]~19 .extended_lut = "off";
defparam \out_data[19]~19 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[19]~19 .shared_arith = "off";

cyclonev_lcell_comb \out_data[20]~20 (
	.dataa(!q_a_20),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[20]~20 .extended_lut = "off";
defparam \out_data[20]~20 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[20]~20 .shared_arith = "off";

cyclonev_lcell_comb \out_data[21]~21 (
	.dataa(!q_a_21),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[21]~21 .extended_lut = "off";
defparam \out_data[21]~21 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \out_data[22]~22 (
	.dataa(!q_a_22),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[22]~22 .extended_lut = "off";
defparam \out_data[22]~22 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[22]~22 .shared_arith = "off";

cyclonev_lcell_comb \out_data[23]~23 (
	.dataa(!q_a_23),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[23]~23 .extended_lut = "off";
defparam \out_data[23]~23 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[23]~23 .shared_arith = "off";

cyclonev_lcell_comb \out_data[24]~24 (
	.dataa(!q_a_24),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[24]~24 .extended_lut = "off";
defparam \out_data[24]~24 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[24]~24 .shared_arith = "off";

cyclonev_lcell_comb \out_data[25]~25 (
	.dataa(!q_a_25),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[25]~25 .extended_lut = "off";
defparam \out_data[25]~25 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[25]~25 .shared_arith = "off";

cyclonev_lcell_comb \out_data[26]~26 (
	.dataa(!q_a_26),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[26]~26 .extended_lut = "off";
defparam \out_data[26]~26 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[26]~26 .shared_arith = "off";

cyclonev_lcell_comb \out_data[27]~27 (
	.dataa(!q_a_27),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[27]~27 .extended_lut = "off";
defparam \out_data[27]~27 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[27]~27 .shared_arith = "off";

cyclonev_lcell_comb \out_data[28]~28 (
	.dataa(!q_a_28),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[28]~28 .extended_lut = "off";
defparam \out_data[28]~28 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[28]~28 .shared_arith = "off";

cyclonev_lcell_comb \out_data[29]~29 (
	.dataa(!q_a_29),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[29]~29 .extended_lut = "off";
defparam \out_data[29]~29 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[29]~29 .shared_arith = "off";

cyclonev_lcell_comb \out_data[30]~30 (
	.dataa(!q_a_30),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[30]~30 .extended_lut = "off";
defparam \out_data[30]~30 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \out_data[31]~31 (
	.dataa(!q_a_31),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem[0][31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[31]~31 .extended_lut = "off";
defparam \out_data[31]~31 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \out_data[31]~31 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!mem_112_0),
	.datab(!mem_used_01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \read~1 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!read_latency_shift_reg_0),
	.datad(!mem_used_0),
	.datae(!src0_valid),
	.dataf(!\read~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~1 .extended_lut = "off";
defparam \read~1 .lut_mask = 64'h0333055500000000;
defparam \read~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!q_a_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(gnd),
	.datad(!mem_used_0),
	.datae(!src0_valid),
	.dataf(!\read~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFF33FF55FF00FF00;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!q_a_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!q_a_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!q_a_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][3]~q ),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!q_a_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][4]~q ),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!q_a_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][5]~q ),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!q_a_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][6]~q ),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!q_a_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][7]~q ),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!q_a_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][8]~q ),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!q_a_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][9]~q ),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!q_a_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][10]~q ),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!q_a_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][11]~q ),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!q_a_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][12]~q ),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!q_a_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][13]~q ),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!q_a_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][14]~q ),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!q_a_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][15]~q ),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!q_a_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][16]~q ),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!q_a_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][17]~q ),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!q_a_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][18]~q ),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!q_a_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][19]~q ),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!q_a_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][20]~q ),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!q_a_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][21]~q ),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!q_a_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][22]~q ),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!q_a_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][23]~q ),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!q_a_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][24]~q ),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!q_a_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][25]~q ),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!q_a_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][26]~q ),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!q_a_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][27]~q ),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!q_a_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][28]~q ),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!q_a_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][29]~q ),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!q_a_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][30]~q ),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!q_a_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][31]~q ),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

endmodule

module soc_system_altera_avalon_sc_fifo_1 (
	clk,
	nxt_out_eop,
	mem_used_1,
	in_ready_hold,
	source0_data_34,
	WideOr0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_112_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	in_data_reg_59,
	m0_write,
	reset,
	nxt_out_eop1,
	out_byte_cnt_reg_2,
	comb,
	WideOr01,
	in_data_reg_60,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	nxt_out_eop;
output 	mem_used_1;
input 	in_ready_hold;
input 	source0_data_34;
input 	WideOr0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_112_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
output 	mem_113_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
input 	last_packet_beat;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
input 	in_data_reg_59;
input 	m0_write;
input 	reset;
input 	nxt_out_eop1;
input 	out_byte_cnt_reg_2;
input 	comb;
input 	WideOr01;
input 	in_data_reg_60;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_88;
input 	in_data_reg_89;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][112]~q ;
wire \mem~0_combout ;
wire \mem~21_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~2_combout ;
wire \mem[1][59]~q ;
wire \mem~1_combout ;
wire \mem[1][60]~q ;
wire \mem~2_combout ;
wire \mem[1][113]~q ;
wire \mem~3_combout ;
wire \mem[1][69]~q ;
wire \mem~4_combout ;
wire \mem[1][68]~q ;
wire \mem~5_combout ;
wire \mem[1][67]~q ;
wire \mem~6_combout ;
wire \mem[1][66]~q ;
wire \mem~7_combout ;
wire \mem[1][65]~q ;
wire \mem~8_combout ;
wire \mem[1][88]~q ;
wire \mem~9_combout ;
wire \mem[1][89]~q ;
wire \mem~10_combout ;
wire \mem[1][90]~q ;
wire \mem~11_combout ;
wire \mem[1][91]~q ;
wire \mem~12_combout ;
wire \mem[1][92]~q ;
wire \mem~13_combout ;
wire \mem[1][93]~q ;
wire \mem~14_combout ;
wire \mem[1][94]~q ;
wire \mem~15_combout ;
wire \mem[1][95]~q ;
wire \mem~16_combout ;
wire \mem[1][96]~q ;
wire \mem~17_combout ;
wire \mem[1][97]~q ;
wire \mem~18_combout ;
wire \mem[1][98]~q ;
wire \mem~19_combout ;
wire \mem[1][99]~q ;
wire \mem~20_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][88] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_88_0),
	.prn(vcc));
defparam \mem[0][88] .is_wysiwyg = "true";
defparam \mem[0][88] .power_up = "low";

dffeas \mem[0][89] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_89_0),
	.prn(vcc));
defparam \mem[0][89] .is_wysiwyg = "true";
defparam \mem[0][89] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!in_ready_hold),
	.datab(!source0_data_34),
	.datac(!WideOr0),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h00D500D500D500D5;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!nxt_out_eop1),
	.datab(!nxt_out_eop),
	.datac(!in_data_reg_59),
	.datad(!in_data_reg_60),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h000007FF000007FF;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!comb),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!WideOr01),
	.dataf(!\write~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h555551550F0F070F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!source0_data_34),
	.datab(!WideOr0),
	.datac(!in_data_reg_60),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h0808080808080808;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem~21 (
	.dataa(!out_valid_reg),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][112]~q ),
	.datad(!nxt_out_eop),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop1),
	.datag(!\mem~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "on";
defparam \mem~21 .lut_mask = 64'h05150F0F15150F0F;
defparam \mem~21 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!comb),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!WideOr01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hCCECCCECCCECCCEC;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!comb),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!WideOr01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h0F0F070F0F0F070F;
defparam \mem_used[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!nxt_out_eop1),
	.datab(!nxt_out_eop),
	.datac(!in_data_reg_59),
	.datad(!in_data_reg_60),
	.datae(!\write~0_combout ),
	.dataf(!\mem_used[0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'h000007FFFFFFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!\mem[1][113]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h2A7F2A7F2A7F2A7F;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h0257025702570257;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][88] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][88]~q ),
	.prn(vcc));
defparam \mem[1][88] .is_wysiwyg = "true";
defparam \mem[1][88] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][88]~q ),
	.datac(!in_data_reg_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][89]~q ),
	.datac(!in_data_reg_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][90]~q ),
	.datac(!in_data_reg_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_axi_master_ni (
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	outclk_wire_0,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	Add45,
	Add55,
	address_burst_6,
	address_burst_7,
	address_burst_8,
	address_burst_9,
	address_burst_10,
	address_burst_11,
	address_burst_12,
	address_burst_13,
	address_burst_14,
	Add56,
	Add46,
	nxt_out_eop,
	new_burst_reg,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	saved_grant_0,
	awready,
	src_valid,
	wready,
	sop_enable1,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	Add1,
	log2ceil,
	src_payload,
	Add3,
	log2ceil1,
	out_data_1,
	log2ceil2,
	src_payload1,
	Add31,
	out_data_0,
	src_payload2,
	out_data_2,
	Selector17,
	out_data_3,
	src_payload3,
	out_data_4,
	src_payload4,
	out_data_5,
	altera_reset_synchronizer_int_chain_out)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	outclk_wire_0;
output 	Add4;
output 	Add5;
output 	Add41;
output 	Add51;
output 	Add42;
output 	Add52;
output 	Add43;
output 	Add53;
output 	Add44;
output 	Add54;
output 	Add45;
output 	Add55;
output 	address_burst_6;
output 	address_burst_7;
output 	address_burst_8;
output 	address_burst_9;
output 	address_burst_10;
output 	address_burst_11;
output 	address_burst_12;
output 	address_burst_13;
output 	address_burst_14;
output 	Add56;
output 	Add46;
input 	nxt_out_eop;
input 	new_burst_reg;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	nxt_in_ready3;
input 	saved_grant_0;
output 	awready;
input 	src_valid;
output 	wready;
output 	sop_enable1;
output 	burst_bytecount_6;
output 	write_cp_data_69;
output 	burst_bytecount_5;
output 	write_cp_data_68;
output 	burst_bytecount_4;
output 	write_cp_data_67;
output 	burst_bytecount_2;
output 	write_cp_data_65;
output 	burst_bytecount_3;
output 	write_cp_data_66;
output 	Add1;
output 	log2ceil;
input 	src_payload;
output 	Add3;
output 	log2ceil1;
output 	out_data_1;
output 	log2ceil2;
input 	src_payload1;
output 	Add31;
output 	out_data_0;
input 	src_payload2;
output 	out_data_2;
output 	Selector17;
output 	out_data_3;
input 	src_payload3;
output 	out_data_4;
input 	src_payload4;
output 	out_data_5;
input 	altera_reset_synchronizer_int_chain_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~7_combout ;
wire \Add4~2 ;
wire \Add5~2 ;
wire \Add4~6 ;
wire \Add5~6 ;
wire \Add4~10 ;
wire \Add5~10 ;
wire \Add4~14 ;
wire \Add5~14 ;
wire \Add4~18 ;
wire \Add5~18 ;
wire \Add4~22 ;
wire \Add5~22 ;
wire \Decoder0~0_combout ;
wire \Decoder1~0_combout ;
wire \Decoder0~1_combout ;
wire \Decoder1~1_combout ;
wire \Decoder0~2_combout ;
wire \Decoder1~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder1~3_combout ;
wire \Decoder0~4_combout ;
wire \Decoder1~4_combout ;
wire \Decoder0~5_combout ;
wire \Decoder1~5_combout ;
wire \Decoder1~6_combout ;
wire \Decoder0~6_combout ;
wire \sop_enable~0_combout ;
wire \Add7~0_combout ;
wire \Add6~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;


soc_system_altera_merlin_address_alignment align_address_to_size(
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.clk(outclk_wire_0),
	.address_burst_6(address_burst_6),
	.address_burst_7(address_burst_7),
	.address_burst_8(address_burst_8),
	.address_burst_9(address_burst_9),
	.address_burst_10(address_burst_10),
	.address_burst_11(address_burst_11),
	.address_burst_12(address_burst_12),
	.address_burst_13(address_burst_13),
	.address_burst_14(address_burst_14),
	.wready(wready),
	.sop_enable(sop_enable1),
	.Add1(Add1),
	.log2ceil(log2ceil),
	.src_payload(src_payload),
	.out_data_1(out_data_1),
	.src_payload1(src_payload1),
	.out_data_0(out_data_0),
	.src_payload2(src_payload2),
	.out_data_2(out_data_2),
	.Selector17(Selector17),
	.out_data_3(out_data_3),
	.src_payload3(src_payload3),
	.out_data_4(out_data_4),
	.src_payload4(src_payload4),
	.out_data_5(out_data_5),
	.reset(altera_reset_synchronizer_int_chain_out),
	.Decoder0(\Decoder0~0_combout ),
	.Decoder01(\Decoder0~1_combout ),
	.Decoder02(\Decoder0~2_combout ),
	.Decoder03(\Decoder0~3_combout ),
	.Decoder04(\Decoder0~4_combout ),
	.Decoder05(\Decoder0~5_combout ),
	.Decoder06(\Decoder0~6_combout ),
	.Decoder07(\Decoder0~7_combout ));

cyclonev_lcell_comb \Decoder0~7 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~7 .extended_lut = "off";
defparam \Decoder0~7 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~7 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add4),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add41),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add42),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add52),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add43),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add53),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add44),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add54),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h00000000000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add45),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h00000000000000FF;
defparam \Add4~21 .shared_arith = "off";

cyclonev_lcell_comb \Add5~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add55),
	.cout(\Add5~22 ),
	.shareout());
defparam \Add5~21 .extended_lut = "off";
defparam \Add5~21 .lut_mask = 64'h00000000000000FF;
defparam \Add5~21 .shared_arith = "off";

cyclonev_lcell_comb \Add5~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add56),
	.cout(),
	.shareout());
defparam \Add5~25 .extended_lut = "off";
defparam \Add5~25 .lut_mask = 64'h00000000000000FF;
defparam \Add5~25 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add46),
	.cout(),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h00000000000000FF;
defparam \Add4~25 .shared_arith = "off";

cyclonev_lcell_comb \awready~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WLAST_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!nxt_in_ready3),
	.datae(!saved_grant_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awready),
	.sumout(),
	.cout(),
	.shareout());
defparam \awready~0 .extended_lut = "off";
defparam \awready~0 .lut_mask = 64'h0000010000000100;
defparam \awready~0 .shared_arith = "off";

cyclonev_lcell_comb \wready~0 (
	.dataa(!new_burst_reg),
	.datab(!nxt_in_ready),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready1),
	.datae(!nxt_in_ready2),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wready),
	.sumout(),
	.cout(),
	.shareout());
defparam \wready~0 .extended_lut = "off";
defparam \wready~0 .lut_mask = 64'h0000000013FFFFFF;
defparam \wready~0 .shared_arith = "off";

dffeas sop_enable(
	.clk(outclk_wire_0),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

dffeas \burst_bytecount[6] (
	.clk(outclk_wire_0),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[69]~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_6),
	.datad(!\Add6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[69]~0 .extended_lut = "off";
defparam \write_cp_data[69]~0 .lut_mask = 64'h0347034703470347;
defparam \write_cp_data[69]~0 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(outclk_wire_0),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[68]~1 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!\Add6~0_combout ),
	.datad(!burst_bytecount_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[68]~1 .extended_lut = "off";
defparam \write_cp_data[68]~1 .lut_mask = 64'h487B487B487B487B;
defparam \write_cp_data[68]~1 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(outclk_wire_0),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[67]~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[67]~2 .extended_lut = "off";
defparam \write_cp_data[67]~2 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[67]~2 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(outclk_wire_0),
	.d(write_cp_data_65),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[65]~3 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_65),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[65]~3 .extended_lut = "off";
defparam \write_cp_data[65]~3 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[65]~3 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(outclk_wire_0),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[66]~4 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[66]~4 .extended_lut = "off";
defparam \write_cp_data[66]~4 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[66]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_lw_AWLEN_1),
	.datab(!h2f_lw_AWLEN_2),
	.datac(!h2f_lw_AWLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~1 (
	.dataa(!h2f_lw_ARLEN_1),
	.datab(!h2f_lw_ARLEN_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil1),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~1 .extended_lut = "off";
defparam \log2ceil~1 .lut_mask = 64'h8888888888888888;
defparam \log2ceil~1 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil2),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~2 .extended_lut = "off";
defparam \log2ceil~2 .lut_mask = 64'h4F004F004F004F00;
defparam \log2ceil~2 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000F003F007F00;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h0808080808080808;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~5 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~5 .extended_lut = "off";
defparam \Decoder1~5 .lut_mask = 64'h0404040404040404;
defparam \Decoder1~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~6 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~6 .extended_lut = "off";
defparam \Decoder1~6 .lut_mask = 64'h0202020202020202;
defparam \Decoder1~6 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h0202020202020202;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_69),
	.datac(!write_cp_data_68),
	.datad(!write_cp_data_67),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h6333333363333333;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add6~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~0 .extended_lut = "off";
defparam \Add6~0 .lut_mask = 64'h0101010101010101;
defparam \Add6~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_68),
	.datac(!write_cp_data_67),
	.datad(!write_cp_data_66),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h6333633363336333;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_67),
	.datac(!write_cp_data_66),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h6363636363636363;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!write_cp_data_65),
	.datab(!write_cp_data_66),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h6666666666666666;
defparam \Add7~3 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_address_alignment (
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	clk,
	address_burst_6,
	address_burst_7,
	address_burst_8,
	address_burst_9,
	address_burst_10,
	address_burst_11,
	address_burst_12,
	address_burst_13,
	address_burst_14,
	wready,
	sop_enable,
	Add1,
	log2ceil,
	src_payload,
	out_data_1,
	src_payload1,
	out_data_0,
	src_payload2,
	out_data_2,
	Selector17,
	out_data_3,
	src_payload3,
	out_data_4,
	src_payload4,
	out_data_5,
	reset,
	Decoder0,
	Decoder01,
	Decoder02,
	Decoder03,
	Decoder04,
	Decoder05,
	Decoder06,
	Decoder07)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	clk;
output 	address_burst_6;
output 	address_burst_7;
output 	address_burst_8;
output 	address_burst_9;
output 	address_burst_10;
output 	address_burst_11;
output 	address_burst_12;
output 	address_burst_13;
output 	address_burst_14;
input 	wready;
input 	sop_enable;
input 	Add1;
input 	log2ceil;
input 	src_payload;
output 	out_data_1;
input 	src_payload1;
output 	out_data_0;
input 	src_payload2;
output 	out_data_2;
output 	Selector17;
output 	out_data_3;
input 	src_payload3;
output 	out_data_4;
input 	src_payload4;
output 	out_data_5;
input 	reset;
input 	Decoder0;
input 	Decoder01;
input 	Decoder02;
input 	Decoder03;
input 	Decoder04;
input 	Decoder05;
input 	Decoder06;
input 	Decoder07;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~5_sumout ;
wire \Add0~5_sumout ;
wire \Selector20~0_combout ;
wire \address_burst[0]~q ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \Selector19~0_combout ;
wire \address_burst[1]~q ;
wire \Add1~2 ;
wire \Add1~9_sumout ;
wire \Add0~2 ;
wire \Add0~9_sumout ;
wire \Selector18~0_combout ;
wire \address_burst[2]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Selector17~1_combout ;
wire \address_burst[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Selector16~0_combout ;
wire \address_burst[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Selector15~0_combout ;
wire \address_burst[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \out_data[6]~6_combout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \out_data[7]~7_combout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \out_data[8]~8_combout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \out_data[9]~9_combout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \out_data[10]~10_combout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \out_data[11]~11_combout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \out_data[12]~12_combout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \out_data[13]~13_combout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \out_data[14]~14_combout ;


dffeas \address_burst[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(\out_data[6]~6_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_6),
	.prn(vcc));
defparam \address_burst[6] .is_wysiwyg = "true";
defparam \address_burst[6] .power_up = "low";

dffeas \address_burst[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(\out_data[7]~7_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_7),
	.prn(vcc));
defparam \address_burst[7] .is_wysiwyg = "true";
defparam \address_burst[7] .power_up = "low";

dffeas \address_burst[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(\out_data[8]~8_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_8),
	.prn(vcc));
defparam \address_burst[8] .is_wysiwyg = "true";
defparam \address_burst[8] .power_up = "low";

dffeas \address_burst[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(\out_data[9]~9_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_9),
	.prn(vcc));
defparam \address_burst[9] .is_wysiwyg = "true";
defparam \address_burst[9] .power_up = "low";

dffeas \address_burst[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(\out_data[10]~10_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_10),
	.prn(vcc));
defparam \address_burst[10] .is_wysiwyg = "true";
defparam \address_burst[10] .power_up = "low";

dffeas \address_burst[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(\out_data[11]~11_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_11),
	.prn(vcc));
defparam \address_burst[11] .is_wysiwyg = "true";
defparam \address_burst[11] .power_up = "low";

dffeas \address_burst[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(\out_data[12]~12_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_12),
	.prn(vcc));
defparam \address_burst[12] .is_wysiwyg = "true";
defparam \address_burst[12] .power_up = "low";

dffeas \address_burst[13] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(\out_data[13]~13_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_13),
	.prn(vcc));
defparam \address_burst[13] .is_wysiwyg = "true";
defparam \address_burst[13] .power_up = "low";

dffeas \address_burst[14] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(\out_data[14]~14_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(wready),
	.q(address_burst_14),
	.prn(vcc));
defparam \address_burst[14] .is_wysiwyg = "true";
defparam \address_burst[14] .power_up = "low";

cyclonev_lcell_comb \out_data[1]~0 (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!sop_enable),
	.datac(!\address_burst[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~0 .extended_lut = "off";
defparam \out_data[1]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~1 (
	.dataa(!h2f_lw_AWADDR_0),
	.datab(!sop_enable),
	.datac(!\address_burst[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~1 .extended_lut = "off";
defparam \out_data[0]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~2 (
	.dataa(!h2f_lw_AWADDR_2),
	.datab(!sop_enable),
	.datac(!\address_burst[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~2 .extended_lut = "off";
defparam \out_data[2]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!Add1),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~3 (
	.dataa(!h2f_lw_AWADDR_3),
	.datab(!sop_enable),
	.datac(!\address_burst[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~3 .extended_lut = "off";
defparam \out_data[3]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~4 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!sop_enable),
	.datac(!\address_burst[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~4 .extended_lut = "off";
defparam \out_data[4]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~5 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!\address_burst[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~5 .extended_lut = "off";
defparam \out_data[5]~5 .lut_mask = 64'h4747474747474747;
defparam \out_data[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[0]~q ),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(!\address_burst[0]~q ),
	.datac(!h2f_lw_AWADDR_0),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!Decoder01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload1),
	.datad(!out_data_0),
	.datae(!\Add1~5_sumout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector20~0 .shared_arith = "off";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[0]~q ),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload),
	.datad(!out_data_1),
	.datae(!\Add1~1_sumout ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector19~0 .shared_arith = "off";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[1]~q ),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload2),
	.datad(!out_data_2),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector18~0 .shared_arith = "off";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[2]~q ),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector17),
	.datad(!out_data_3),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~1 .extended_lut = "off";
defparam \Selector17~1 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector17~1 .shared_arith = "off";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector17~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[3]~q ),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload3),
	.datad(!out_data_4),
	.datae(!\Add1~17_sumout ),
	.dataf(!\Add0~17_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector16~0 .shared_arith = "off";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[4]~q ),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_5),
	.datad(!Decoder05),
	.datae(gnd),
	.dataf(!\address_burst[5]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_5),
	.datad(!Decoder05),
	.datae(gnd),
	.dataf(!\address_burst[5]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload4),
	.datad(!out_data_5),
	.datae(!\Add1~21_sumout ),
	.dataf(!\Add0~21_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector15~0 .shared_arith = "off";

dffeas \address_burst[5] (
	.clk(clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[5]~q ),
	.prn(vcc));
defparam \address_burst[5] .is_wysiwyg = "true";
defparam \address_burst[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_6),
	.datad(!Decoder06),
	.datae(gnd),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~6 (
	.dataa(!h2f_lw_AWADDR_6),
	.datab(!sop_enable),
	.datac(!address_burst_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~6 .extended_lut = "off";
defparam \out_data[6]~6 .lut_mask = 64'h4747474747474747;
defparam \out_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_7),
	.datad(!Decoder07),
	.datae(gnd),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~7 (
	.dataa(!h2f_lw_AWADDR_7),
	.datab(!sop_enable),
	.datac(!address_burst_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~7 .extended_lut = "off";
defparam \out_data[7]~7 .lut_mask = 64'h4747474747474747;
defparam \out_data[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_8),
	.datad(!address_burst_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~8 (
	.dataa(!h2f_lw_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~8 .extended_lut = "off";
defparam \out_data[8]~8 .lut_mask = 64'h4747474747474747;
defparam \out_data[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_9),
	.datad(!address_burst_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~9 (
	.dataa(!h2f_lw_AWADDR_9),
	.datab(!sop_enable),
	.datac(!address_burst_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~9 .extended_lut = "off";
defparam \out_data[9]~9 .lut_mask = 64'h4747474747474747;
defparam \out_data[9]~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_10),
	.datad(!address_burst_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~10 (
	.dataa(!h2f_lw_AWADDR_10),
	.datab(!sop_enable),
	.datac(!address_burst_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~10 .extended_lut = "off";
defparam \out_data[10]~10 .lut_mask = 64'h4747474747474747;
defparam \out_data[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_11),
	.datad(!address_burst_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~11 (
	.dataa(!h2f_lw_AWADDR_11),
	.datab(!sop_enable),
	.datac(!address_burst_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~11 .extended_lut = "off";
defparam \out_data[11]~11 .lut_mask = 64'h4747474747474747;
defparam \out_data[11]~11 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_12),
	.datad(!address_burst_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~12 (
	.dataa(!h2f_lw_AWADDR_12),
	.datab(!sop_enable),
	.datac(!address_burst_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~12 .extended_lut = "off";
defparam \out_data[12]~12 .lut_mask = 64'h4747474747474747;
defparam \out_data[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_13),
	.datad(!address_burst_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~13 (
	.dataa(!h2f_lw_AWADDR_13),
	.datab(!sop_enable),
	.datac(!address_burst_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~13 .extended_lut = "off";
defparam \out_data[13]~13 .lut_mask = 64'h4747474747474747;
defparam \out_data[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_14),
	.datad(!address_burst_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~14 (
	.dataa(!h2f_lw_AWADDR_14),
	.datab(!sop_enable),
	.datac(!address_burst_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~14 .extended_lut = "off";
defparam \out_data[14]~14 .lut_mask = 64'h4747474747474747;
defparam \out_data[14]~14 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_burst_adapter (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	outclk_wire_0,
	address_burst_6,
	address_burst_7,
	address_burst_8,
	address_burst_9,
	address_burst_10,
	address_burst_11,
	address_burst_12,
	address_burst_13,
	address_burst_14,
	nxt_out_eop,
	saved_grant_1,
	new_burst_reg,
	mem_used_1,
	in_ready_hold,
	in_narrow_reg,
	source0_data_33,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	source0_data_35,
	in_byteen_reg_3,
	source0_data_351,
	in_byteen_reg_1,
	source0_data_331,
	WideOr0,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	saved_grant_0,
	src_valid,
	in_data_reg_59,
	in_data_reg_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	int_nxt_addr_reg_dly_10,
	int_nxt_addr_reg_dly_11,
	int_nxt_addr_reg_dly_12,
	int_nxt_addr_reg_dly_13,
	int_nxt_addr_reg_dly_14,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	source0_data_332,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	source0_data_352,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	altera_reset_synchronizer_int_chain_out,
	WideOr1,
	src_payload_0,
	nxt_out_eop1,
	out_byte_cnt_reg_2,
	sop_enable,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_77,
	src_payload,
	src_data_71,
	out_data_1,
	src_payload1,
	src_data_70,
	out_data_0,
	src_data_34,
	src_data_32,
	src_data_35,
	src_data_33,
	cp_ready,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	src_payload2,
	src_payload3,
	src_data_72,
	out_data_2,
	src_payload4,
	src_data_73,
	out_data_3,
	src_payload5,
	src_data_74,
	out_data_4,
	src_payload6,
	src_data_75,
	out_data_5,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_data_711,
	src_data_701,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_721,
	src_data_731,
	src_data_741,
	src_data_751,
	src_data_76,
	src_data_761,
	src_data_762)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARADDR_6;
input 	h2f_lw_ARADDR_7;
input 	h2f_lw_ARADDR_8;
input 	h2f_lw_ARADDR_9;
input 	h2f_lw_ARADDR_10;
input 	h2f_lw_ARADDR_11;
input 	h2f_lw_ARADDR_12;
input 	h2f_lw_ARADDR_13;
input 	h2f_lw_ARADDR_14;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	outclk_wire_0;
input 	address_burst_6;
input 	address_burst_7;
input 	address_burst_8;
input 	address_burst_9;
input 	address_burst_10;
input 	address_burst_11;
input 	address_burst_12;
input 	address_burst_13;
input 	address_burst_14;
output 	nxt_out_eop;
input 	saved_grant_1;
output 	new_burst_reg;
input 	mem_used_1;
output 	in_ready_hold;
output 	in_narrow_reg;
output 	source0_data_33;
output 	in_byteen_reg_2;
output 	source0_data_34;
output 	in_byteen_reg_0;
output 	source0_data_32;
output 	source0_data_35;
output 	in_byteen_reg_3;
output 	source0_data_351;
output 	in_byteen_reg_1;
output 	source0_data_331;
input 	WideOr0;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
output 	nxt_in_ready3;
input 	saved_grant_0;
input 	src_valid;
output 	in_data_reg_59;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
output 	int_nxt_addr_reg_dly_10;
output 	int_nxt_addr_reg_dly_11;
output 	int_nxt_addr_reg_dly_12;
output 	int_nxt_addr_reg_dly_13;
output 	int_nxt_addr_reg_dly_14;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	source0_data_332;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	source0_data_352;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	altera_reset_synchronizer_int_chain_out;
input 	WideOr1;
input 	src_payload_0;
output 	nxt_out_eop1;
output 	out_byte_cnt_reg_2;
input 	sop_enable;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_3;
input 	write_cp_data_66;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_77;
input 	src_payload;
input 	src_data_71;
input 	out_data_1;
input 	src_payload1;
input 	src_data_70;
input 	out_data_0;
input 	src_data_34;
input 	src_data_32;
input 	src_data_35;
input 	src_data_33;
input 	cp_ready;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
input 	src_payload2;
input 	src_payload3;
input 	src_data_72;
input 	out_data_2;
input 	src_payload4;
input 	src_data_73;
input 	out_data_3;
input 	src_payload5;
input 	src_data_74;
input 	out_data_4;
input 	src_payload6;
input 	src_data_75;
input 	out_data_5;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_data_711;
input 	src_data_701;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_721;
input 	src_data_731;
input 	src_data_741;
input 	src_data_751;
input 	src_data_76;
input 	src_data_761;
input 	src_data_762;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARADDR_5(h2f_lw_ARADDR_5),
	.h2f_lw_ARADDR_6(h2f_lw_ARADDR_6),
	.h2f_lw_ARADDR_7(h2f_lw_ARADDR_7),
	.h2f_lw_ARADDR_8(h2f_lw_ARADDR_8),
	.h2f_lw_ARADDR_9(h2f_lw_ARADDR_9),
	.h2f_lw_ARADDR_10(h2f_lw_ARADDR_10),
	.h2f_lw_ARADDR_11(h2f_lw_ARADDR_11),
	.h2f_lw_ARADDR_12(h2f_lw_ARADDR_12),
	.h2f_lw_ARADDR_13(h2f_lw_ARADDR_13),
	.h2f_lw_ARADDR_14(h2f_lw_ARADDR_14),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.outclk_wire_0(outclk_wire_0),
	.address_burst_6(address_burst_6),
	.address_burst_7(address_burst_7),
	.address_burst_8(address_burst_8),
	.address_burst_9(address_burst_9),
	.address_burst_10(address_burst_10),
	.address_burst_11(address_burst_11),
	.address_burst_12(address_burst_12),
	.address_burst_13(address_burst_13),
	.address_burst_14(address_burst_14),
	.nxt_out_eop(nxt_out_eop),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,src_data_762,src_data_751,
src_data_741,src_data_731,src_data_721,src_data_711,src_data_701,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload37,src_payload36,
src_payload35,src_payload34,src_payload33,src_payload32,src_payload31,src_payload30,src_payload29,src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,
src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload2}),
	.new_burst_reg1(new_burst_reg),
	.mem_used_1(mem_used_1),
	.in_ready_hold1(in_ready_hold),
	.in_narrow_reg1(in_narrow_reg),
	.source0_data_33(source0_data_33),
	.in_byteen_reg_2(in_byteen_reg_2),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(in_byteen_reg_0),
	.source0_data_32(source0_data_32),
	.source0_data_35(source0_data_35),
	.in_byteen_reg_3(in_byteen_reg_3),
	.source0_data_351(source0_data_351),
	.in_byteen_reg_1(in_byteen_reg_1),
	.source0_data_331(source0_data_331),
	.WideOr0(WideOr0),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.nxt_in_ready2(nxt_in_ready2),
	.nxt_in_ready3(nxt_in_ready3),
	.src_valid(src_valid),
	.in_data_reg_59(in_data_reg_59),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_5(int_nxt_addr_reg_dly_5),
	.int_nxt_addr_reg_dly_6(int_nxt_addr_reg_dly_6),
	.int_nxt_addr_reg_dly_7(int_nxt_addr_reg_dly_7),
	.int_nxt_addr_reg_dly_8(int_nxt_addr_reg_dly_8),
	.int_nxt_addr_reg_dly_9(int_nxt_addr_reg_dly_9),
	.int_nxt_addr_reg_dly_10(int_nxt_addr_reg_dly_10),
	.int_nxt_addr_reg_dly_11(int_nxt_addr_reg_dly_11),
	.int_nxt_addr_reg_dly_12(int_nxt_addr_reg_dly_12),
	.int_nxt_addr_reg_dly_13(int_nxt_addr_reg_dly_13),
	.int_nxt_addr_reg_dly_14(int_nxt_addr_reg_dly_14),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.source0_data_332(source0_data_332),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.source0_data_352(source0_data_352),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.WideOr1(WideOr1),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop1(nxt_out_eop1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.sop_enable(sop_enable),
	.burst_bytecount_6(burst_bytecount_6),
	.write_cp_data_69(write_cp_data_69),
	.burst_bytecount_5(burst_bytecount_5),
	.write_cp_data_68(write_cp_data_68),
	.burst_bytecount_4(burst_bytecount_4),
	.write_cp_data_67(write_cp_data_67),
	.burst_bytecount_2(burst_bytecount_2),
	.write_cp_data_65(write_cp_data_65),
	.burst_bytecount_3(burst_bytecount_3),
	.write_cp_data_66(write_cp_data_66),
	.in_data_reg_60(in_data_reg_60),
	.src_payload(src_payload),
	.src_data_71(src_data_71),
	.out_data_1(out_data_1),
	.src_payload1(src_payload1),
	.src_data_70(src_data_70),
	.out_data_0(out_data_0),
	.cp_ready(cp_ready),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_88(in_data_reg_88),
	.in_data_reg_89(in_data_reg_89),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.src_payload2(src_payload3),
	.src_data_72(src_data_72),
	.out_data_2(out_data_2),
	.src_payload3(src_payload4),
	.src_data_73(src_data_73),
	.out_data_3(out_data_3),
	.src_payload4(src_payload5),
	.src_data_74(src_data_74),
	.out_data_4(out_data_4),
	.src_payload5(src_payload6),
	.src_data_75(src_data_75),
	.out_data_5(out_data_5),
	.src_data_76(src_data_76),
	.src_data_761(src_data_761));

endmodule

module soc_system_altera_merlin_burst_adapter_13_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	outclk_wire_0,
	address_burst_6,
	address_burst_7,
	address_burst_8,
	address_burst_9,
	address_burst_10,
	address_burst_11,
	address_burst_12,
	address_burst_13,
	address_burst_14,
	nxt_out_eop,
	sink0_data,
	new_burst_reg1,
	mem_used_1,
	in_ready_hold1,
	in_narrow_reg1,
	source0_data_33,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	source0_data_35,
	in_byteen_reg_3,
	source0_data_351,
	in_byteen_reg_1,
	source0_data_331,
	WideOr0,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	src_valid,
	in_data_reg_59,
	in_data_reg_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	int_nxt_addr_reg_dly_10,
	int_nxt_addr_reg_dly_11,
	int_nxt_addr_reg_dly_12,
	int_nxt_addr_reg_dly_13,
	int_nxt_addr_reg_dly_14,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	source0_data_332,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	source0_data_352,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	altera_reset_synchronizer_int_chain_out,
	WideOr1,
	sink0_endofpacket,
	nxt_out_eop1,
	out_byte_cnt_reg_2,
	sop_enable,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_3,
	write_cp_data_66,
	in_data_reg_60,
	src_payload,
	src_data_71,
	out_data_1,
	src_payload1,
	src_data_70,
	out_data_0,
	cp_ready,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	src_payload2,
	src_data_72,
	out_data_2,
	src_payload3,
	src_data_73,
	out_data_3,
	src_payload4,
	src_data_74,
	out_data_4,
	src_payload5,
	src_data_75,
	out_data_5,
	src_data_76,
	src_data_761)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARADDR_6;
input 	h2f_lw_ARADDR_7;
input 	h2f_lw_ARADDR_8;
input 	h2f_lw_ARADDR_9;
input 	h2f_lw_ARADDR_10;
input 	h2f_lw_ARADDR_11;
input 	h2f_lw_ARADDR_12;
input 	h2f_lw_ARADDR_13;
input 	h2f_lw_ARADDR_14;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	outclk_wire_0;
input 	address_burst_6;
input 	address_burst_7;
input 	address_burst_8;
input 	address_burst_9;
input 	address_burst_10;
input 	address_burst_11;
input 	address_burst_12;
input 	address_burst_13;
input 	address_burst_14;
output 	nxt_out_eop;
input 	[111:0] sink0_data;
output 	new_burst_reg1;
input 	mem_used_1;
output 	in_ready_hold1;
output 	in_narrow_reg1;
output 	source0_data_33;
output 	in_byteen_reg_2;
output 	source0_data_34;
output 	in_byteen_reg_0;
output 	source0_data_32;
output 	source0_data_35;
output 	in_byteen_reg_3;
output 	source0_data_351;
output 	in_byteen_reg_1;
output 	source0_data_331;
input 	WideOr0;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
output 	nxt_in_ready3;
input 	src_valid;
output 	in_data_reg_59;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
output 	int_nxt_addr_reg_dly_10;
output 	int_nxt_addr_reg_dly_11;
output 	int_nxt_addr_reg_dly_12;
output 	int_nxt_addr_reg_dly_13;
output 	int_nxt_addr_reg_dly_14;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	source0_data_332;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	source0_data_352;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	altera_reset_synchronizer_int_chain_out;
input 	WideOr1;
input 	sink0_endofpacket;
output 	nxt_out_eop1;
output 	out_byte_cnt_reg_2;
input 	sop_enable;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_3;
input 	write_cp_data_66;
output 	in_data_reg_60;
input 	src_payload;
input 	src_data_71;
input 	out_data_1;
input 	src_payload1;
input 	src_data_70;
input 	out_data_0;
input 	cp_ready;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
input 	src_payload2;
input 	src_data_72;
input 	out_data_2;
input 	src_payload3;
input 	src_data_73;
input 	out_data_3;
input 	src_payload4;
input 	src_data_74;
input 	out_data_4;
input 	src_payload5;
input 	src_data_75;
input 	out_data_5;
input 	src_data_76;
input 	src_data_761;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \WideNor0~0_combout ;
wire \WideNor0~1_combout ;
wire \in_valid~combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~3_combout ;
wire \Selector1~0_combout ;
wire \Selector1~4_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~3_combout ;
wire \Selector3~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \WideOr0~0_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \nxt_in_ready~5_combout ;
wire \Selector1~5_combout ;
wire \Selector1~6_combout ;
wire \state.ST_COMP_TRANS~q ;
wire \in_eop_reg~q ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \d0_int_bytes_remaining[2]~8_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~7_combout ;
wire \d0_int_bytes_remaining[3]~9_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~2_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \d0_int_bytes_remaining[4]~5_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \Selector1~2_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \LessThan0~0_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \d0_in_size[0]~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \d0_int_nxt_addr[0]~4_combout ;
wire \d0_int_nxt_addr[0]~5_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~0_combout ;
wire \d0_int_nxt_addr[1]~1_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \source0_data[34]~1_combout ;
wire \nxt_out_valid~0_combout ;
wire \Selector3~1_combout ;
wire \nxt_in_ready~2_combout ;
wire \d0_in_size[2]~1_combout ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \Add0~2 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~6_combout ;
wire \d0_int_nxt_addr[2]~7_combout ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~8_combout ;
wire \d0_int_nxt_addr[3]~9_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[4]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \in_burstwrap_reg[4]~q ;
wire \nxt_addr[4]~combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \d0_int_nxt_addr[4]~10_combout ;
wire \d0_int_nxt_addr[4]~11_combout ;
wire \ShiftLeft0~5_combout ;
wire \int_byte_cnt_narrow_reg[5]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \in_burstwrap_reg[5]~q ;
wire \nxt_addr[5]~combout ;
wire \int_nxt_addr_reg[5]~q ;
wire \d0_int_nxt_addr[5]~12_combout ;
wire \d0_int_nxt_addr[5]~13_combout ;
wire \d0_int_nxt_addr[6]~14_combout ;
wire \in_burstwrap_reg[6]~q ;
wire \nxt_addr[6]~8_combout ;
wire \int_nxt_addr_reg[6]~q ;
wire \ShiftLeft0~6_combout ;
wire \int_byte_cnt_narrow_reg[6]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \d0_int_nxt_addr[6]~15_combout ;
wire \d0_int_nxt_addr[7]~16_combout ;
wire \nxt_addr[7]~7_combout ;
wire \int_nxt_addr_reg[7]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \d0_int_nxt_addr[7]~17_combout ;
wire \d0_int_nxt_addr[8]~18_combout ;
wire \nxt_addr[8]~6_combout ;
wire \int_nxt_addr_reg[8]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \d0_int_nxt_addr[8]~19_combout ;
wire \d0_int_nxt_addr[9]~20_combout ;
wire \nxt_addr[9]~5_combout ;
wire \int_nxt_addr_reg[9]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \d0_int_nxt_addr[9]~21_combout ;
wire \d0_int_nxt_addr[10]~22_combout ;
wire \nxt_addr[10]~4_combout ;
wire \int_nxt_addr_reg[10]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \d0_int_nxt_addr[10]~23_combout ;
wire \d0_int_nxt_addr[11]~24_combout ;
wire \nxt_addr[11]~3_combout ;
wire \int_nxt_addr_reg[11]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \d0_int_nxt_addr[11]~25_combout ;
wire \d0_int_nxt_addr[12]~26_combout ;
wire \nxt_addr[12]~2_combout ;
wire \int_nxt_addr_reg[12]~q ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \d0_int_nxt_addr[12]~27_combout ;
wire \d0_int_nxt_addr[13]~28_combout ;
wire \nxt_addr[13]~1_combout ;
wire \int_nxt_addr_reg[13]~q ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \d0_int_nxt_addr[13]~29_combout ;
wire \d0_int_nxt_addr[14]~30_combout ;
wire \nxt_addr[14]~0_combout ;
wire \int_nxt_addr_reg[14]~q ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \d0_int_nxt_addr[14]~31_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~5_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~6_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~7_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~8_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~9_combout ;


soc_system_altera_merlin_address_alignment_1 align_address_to_size(
	.ShiftLeft0(\ShiftLeft0~0_combout ),
	.d0_in_size_0(\d0_in_size[0]~0_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_out_eop~1 (
	.dataa(!\in_bytecount_reg_zero~q ),
	.datab(!source0_data_34),
	.datac(!WideOr0),
	.datad(!in_ready_hold1),
	.datae(!\state.ST_COMP_TRANS~q ),
	.dataf(!mem_used_1),
	.datag(!\in_eop_reg~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~1 .extended_lut = "on";
defparam \nxt_out_eop~1 .lut_mask = 64'h0F0F15000F0F5555;
defparam \nxt_out_eop~1 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(new_burst_reg1),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

dffeas in_ready_hold(
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

dffeas in_narrow_reg(
	.clk(outclk_wire_0),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \source0_data[33]~0 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_narrow_reg1),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(!\int_nxt_addr_reg_dly[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[33]~0 .extended_lut = "off";
defparam \source0_data[33]~0 .lut_mask = 64'h0111111100000000;
defparam \source0_data[33]~0 .shared_arith = "off";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

cyclonev_lcell_comb \source0_data[34]~2 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_narrow_reg1),
	.datac(!source0_data_33),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(!in_byteen_reg_2),
	.dataf(!\source0_data[34]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[34]~2 .extended_lut = "off";
defparam \source0_data[34]~2 .lut_mask = 64'h110FFFEF000FEEEF;
defparam \source0_data[34]~2 .shared_arith = "off";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

cyclonev_lcell_comb \source0_data[32]~3 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_narrow_reg1),
	.datac(!\int_nxt_addr_reg_dly[1]~q ),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(!in_byteen_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[32]~3 .extended_lut = "off";
defparam \source0_data[32]~3 .lut_mask = 64'h1000FEEE1000FEEE;
defparam \source0_data[32]~3 .shared_arith = "off";

cyclonev_lcell_comb \source0_data[35]~4 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_narrow_reg1),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(!\int_nxt_addr_reg_dly[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~4 .extended_lut = "off";
defparam \source0_data[35]~4 .lut_mask = 64'h0001001100010011;
defparam \source0_data[35]~4 .shared_arith = "off";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

cyclonev_lcell_comb \source0_data[35]~5 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_narrow_reg1),
	.datac(!\in_size_reg[2]~q ),
	.datad(!\in_size_reg[1]~q ),
	.datae(!in_byteen_reg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_351),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~5 .extended_lut = "off";
defparam \source0_data[35]~5 .lut_mask = 64'hFEEE1000FEEE1000;
defparam \source0_data[35]~5 .shared_arith = "off";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

cyclonev_lcell_comb \source0_data[33]~6 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_byteen_reg_1),
	.datac(!in_narrow_reg1),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(!\int_nxt_addr_reg_dly[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_331),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[33]~6 .extended_lut = "off";
defparam \source0_data[33]~6 .lut_mask = 64'h3232373232323732;
defparam \source0_data[33]~6 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!mem_used_1),
	.datac(!in_ready_hold1),
	.datad(!source0_data_34),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h4404040444040404;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_ready_hold1),
	.datac(!out_valid_reg1),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h7250505072505050;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~3 (
	.dataa(!mem_used_1),
	.datab(!in_ready_hold1),
	.datac(!source0_data_34),
	.datad(!WideOr0),
	.datae(!out_valid_reg1),
	.dataf(!\nxt_in_ready~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~3 .extended_lut = "off";
defparam \nxt_in_ready~3 .lut_mask = 64'h00000000FFFFA222;
defparam \nxt_in_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~4 (
	.dataa(!new_burst_reg1),
	.datab(!nxt_in_ready),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready1),
	.datae(!nxt_in_ready2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~4 .extended_lut = "off";
defparam \nxt_in_ready~4 .lut_mask = 64'hEC000000EC000000;
defparam \nxt_in_ready~4 .shared_arith = "off";

dffeas \in_data_reg[59] (
	.clk(outclk_wire_0),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[2]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[3]~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[4]~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[5] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[5]~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_5),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[5] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[5] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[6] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[6]~15_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_6),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[6] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[6] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[7] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[7]~17_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_7),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[7] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[7] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[8] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[8]~19_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_8),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[8] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[8] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[9] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[9]~21_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_9),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[9] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[9] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[10] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[10]~23_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_10),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[10] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[10] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[11] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[11]~25_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_11),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[11] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[11] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[12] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[12]~27_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_12),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[12] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[12] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[13] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[13]~29_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_13),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[13] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[13] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[14] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[14]~31_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_14),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[14] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[14] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

cyclonev_lcell_comb \source0_data[33]~7 (
	.dataa(!source0_data_33),
	.datab(!source0_data_331),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_332),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[33]~7 .extended_lut = "off";
defparam \source0_data[33]~7 .lut_mask = 64'h7777777777777777;
defparam \source0_data[33]~7 .shared_arith = "off";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

cyclonev_lcell_comb \source0_data[35]~8 (
	.dataa(!source0_data_35),
	.datab(!source0_data_351),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_352),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~8 .extended_lut = "off";
defparam \source0_data[35]~8 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \source0_data[35]~8 .shared_arith = "off";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!new_burst_reg1),
	.datac(!mem_used_1),
	.datad(!in_ready_hold1),
	.datae(!source0_data_34),
	.dataf(!WideOr0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h1010001000100010;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \in_data_reg[60] (
	.clk(outclk_wire_0),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[88] (
	.clk(outclk_wire_0),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_88),
	.prn(vcc));
defparam \in_data_reg[88] .is_wysiwyg = "true";
defparam \in_data_reg[88] .power_up = "low";

dffeas \in_data_reg[89] (
	.clk(outclk_wire_0),
	.d(sink0_data[89]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_89),
	.prn(vcc));
defparam \in_data_reg[89] .is_wysiwyg = "true";
defparam \in_data_reg[89] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(outclk_wire_0),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(outclk_wire_0),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(outclk_wire_0),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(outclk_wire_0),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(outclk_wire_0),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(outclk_wire_0),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(outclk_wire_0),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(outclk_wire_0),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sop_enable),
	.datab(!burst_bytecount_6),
	.datac(!burst_bytecount_5),
	.datad(!burst_bytecount_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h4000400040004000;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~1 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!burst_bytecount_2),
	.datad(!burst_bytecount_3),
	.datae(!\WideNor0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~1 .extended_lut = "off";
defparam \WideNor0~1 .lut_mask = 64'h8888A8888888A888;
defparam \WideNor0~1 .shared_arith = "off";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold1),
	.datab(!WideOr1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h1111111111111111;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!new_burst_reg1),
	.datab(!nxt_in_ready),
	.datac(!nxt_out_eop),
	.datad(!nxt_in_ready1),
	.datae(!nxt_in_ready2),
	.dataf(!\in_valid~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0000000013FFFFFF;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(outclk_wire_0),
	.d(\WideNor0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[59]),
	.datae(!\in_valid~combout ),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h000055FFC0C0FFFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!in_ready_hold1),
	.datac(!source0_data_34),
	.datad(!WideOr0),
	.datae(!out_valid_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hFFFFA222FFFFA222;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!sink0_data[60]),
	.datab(!\in_valid~combout ),
	.datac(!\state.ST_IDLE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h1010101010101010;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h2222222222222222;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!\in_valid~combout ),
	.datab(!\Selector1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'h4444444444444444;
defparam \Selector1~4 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!mem_used_1),
	.datab(!in_ready_hold1),
	.datac(!source0_data_34),
	.datad(!WideOr0),
	.datae(!out_valid_reg1),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0000A22200000000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_5),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~0 .lut_mask = 64'h2222822222228222;
defparam \nxt_uncomp_subburst_byte_cnt[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~1 (
	.dataa(!mem_used_1),
	.datab(!in_ready_hold1),
	.datac(!source0_data_34),
	.datad(!WideOr0),
	.datae(!out_valid_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~1 .lut_mask = 64'h0000A2220000A222;
defparam \nxt_uncomp_subburst_byte_cnt~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h0544054405440544;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.datad(!out_uncomp_byte_cnt_reg_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .lut_mask = 64'h0454045404540454;
defparam \nxt_uncomp_subburst_byte_cnt[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop1),
	.datab(!nxt_out_eop),
	.datac(!\nxt_in_ready~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_5),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h00008000AAAA2AAA;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF00011110000B111;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~0_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.datad(!\Selector3~0_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.dataf(!\WideOr0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0000000000800000;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000EAC00000EAC0;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!in_ready_hold1),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!WideOr1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h0000001500000015;
defparam \Selector2~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~3 (
	.dataa(!sink0_data[60]),
	.datab(!in_ready_hold1),
	.datac(!src_valid),
	.datad(!\Selector2~0_combout ),
	.datae(!\Selector2~1_combout ),
	.dataf(!\Selector2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~3 .extended_lut = "off";
defparam \Selector2~3 .lut_mask = 64'h02FF00FFAAFFAAFF;
defparam \Selector2~3 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~5 .extended_lut = "off";
defparam \nxt_in_ready~5 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~5 (
	.dataa(!sink0_data[60]),
	.datab(!\nxt_in_ready~5_combout ),
	.datac(!\in_valid~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~5 .extended_lut = "off";
defparam \Selector1~5 .lut_mask = 64'h0404040404040404;
defparam \Selector1~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~6 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!\Selector1~3_combout ),
	.datae(!\Selector1~4_combout ),
	.dataf(!\Selector1~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~6 .extended_lut = "off";
defparam \Selector1~6 .lut_mask = 64'h40FF55FF7FFF7FFF;
defparam \Selector1~6 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector1~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_COMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!in_ready_hold1),
	.datac(!nxt_out_eop1),
	.datad(!nxt_out_eop),
	.datae(!WideOr1),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h5000511150005000;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~8 (
	.dataa(!new_burst_reg1),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~8 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~7 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~9 (
	.dataa(!new_burst_reg1),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(!\d0_int_bytes_remaining[3]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~9 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~9 .lut_mask = 64'h208A75DF208A75DF;
defparam \d0_int_bytes_remaining[3]~9 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[3]~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'hB4F0B4F0B4F0B4F0;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!sink0_data[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'h001E001E001E001E;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~5 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[59]),
	.datac(!\Add1~2_combout ),
	.datad(!write_cp_data_67),
	.datae(!\d0_int_bytes_remaining[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~5 .lut_mask = 64'hA0B1F5F5A0B1F5F5;
defparam \d0_int_bytes_remaining[4]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[4]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(!\int_bytes_remaining_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hB4F0F0F0B4F0F0F0;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!sink0_data[60]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h000001FE000001FE;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[59]),
	.datac(!\Add1~1_combout ),
	.datad(!write_cp_data_68),
	.datae(!\d0_int_bytes_remaining[5]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'hA0B1F5F5A0B1F5F5;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(!\int_bytes_remaining_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000000040000000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!sink0_data[60]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h0000000100000001;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[59]),
	.datac(!\int_bytes_remaining_reg[6]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!write_cp_data_69),
	.dataf(!\d0_int_bytes_remaining[6]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h0AA01BB15FF55FF5;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop1),
	.datac(!nxt_out_eop),
	.datad(!\nxt_in_ready~5_combout ),
	.datae(!\in_valid~combout ),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h0000555500001500;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!new_burst_reg1),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~6_combout ),
	.datae(!\int_bytes_remaining_reg[3]~q ),
	.dataf(!\d0_int_bytes_remaining[3]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h085D207508082020;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[6]~1_combout ),
	.datac(!\d0_int_bytes_remaining[5]~3_combout ),
	.datad(!\d0_int_bytes_remaining[4]~5_combout ),
	.datae(!\Selector1~2_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAA0000EAAAC000;
defparam \new_burst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[2]~q ),
	.datac(!\in_size_reg[1]~q ),
	.datad(!sink0_data[78]),
	.datae(!sink0_data[79]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'hD5808080D5808080;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_in_size[0]~0 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[0]~q ),
	.datac(!sink0_data[77]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_in_size[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_in_size[0]~0 .extended_lut = "off";
defparam \d0_in_size[0]~0 .lut_mask = 64'h2727272727272727;
defparam \d0_in_size[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\ShiftLeft0~0_combout ),
	.datab(!\d0_in_size[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h1111111111111111;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload1),
	.datad(!src_data_70),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~4 (
	.dataa(!new_burst_reg1),
	.datab(!\ShiftLeft0~0_combout ),
	.datac(!\int_nxt_addr_reg[0]~q ),
	.datad(!\d0_in_size[0]~0_combout ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~4 .lut_mask = 64'h0A0A1B0A0A0A1B0A;
defparam \d0_int_nxt_addr[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~5 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(!\d0_int_nxt_addr[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~5 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[0]~5 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload),
	.datad(!src_data_71),
	.datae(!\in_burstwrap_reg[1]~q ),
	.dataf(!\d0_int_nxt_addr[1]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~0 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~1 (
	.dataa(!new_burst_reg1),
	.datab(!\int_nxt_addr_reg[1]~q ),
	.datac(!\d0_int_nxt_addr[1]~0_combout ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~1 .lut_mask = 64'h2227222722272227;
defparam \d0_int_nxt_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[1]~q ),
	.dataf(!\d0_int_nxt_addr[1]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \source0_data[34]~1 (
	.dataa(!\in_size_reg[2]~q ),
	.datab(!\in_size_reg[1]~q ),
	.datac(!\int_nxt_addr_reg_dly[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source0_data[34]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[34]~1 .extended_lut = "off";
defparam \source0_data[34]~1 .lut_mask = 64'h8080808080808080;
defparam \source0_data[34]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!new_burst_reg1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~0_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.datad(!\Selector3~0_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.dataf(!\WideOr0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h00FF00FF007F00FF;
defparam \Selector3~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!\state.ST_COMP_TRANS~q ),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_in_size[2]~1 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[2]~q ),
	.datac(!sink0_data[79]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_in_size[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_in_size[2]~1 .extended_lut = "off";
defparam \d0_in_size[2]~1 .lut_mask = 64'h2727272727272727;
defparam \d0_in_size[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[1]~q ),
	.datac(!sink0_data[78]),
	.datad(!\d0_in_size[2]~1_combout ),
	.datae(!\d0_in_size[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h2700000027000000;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload2),
	.datad(!src_data_72),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~6 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[59]),
	.datae(!\int_nxt_addr_reg[2]~q ),
	.dataf(!out_data_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~6 .lut_mask = 64'h0101F1F1010FF1FF;
defparam \d0_int_nxt_addr[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~7 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~7 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[1]~q ),
	.datac(!sink0_data[78]),
	.datad(!\d0_in_size[2]~1_combout ),
	.datae(!\d0_in_size[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h0000270000002700;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload3),
	.datad(!src_data_73),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~8 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[59]),
	.datae(!\int_nxt_addr_reg[3]~q ),
	.dataf(!out_data_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~8 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~8 .lut_mask = 64'h0101F1F1010FF1FF;
defparam \d0_int_nxt_addr[3]~8 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~9 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~9 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~9 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[3]~9 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[1]~q ),
	.datac(!sink0_data[78]),
	.datad(!\d0_in_size[2]~1_combout ),
	.datae(!\d0_in_size[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h00D8000000D80000;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[4] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[4]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[4] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[4]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[74]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[4] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload4),
	.datad(!src_data_74),
	.datae(!\in_burstwrap_reg[4]~q ),
	.dataf(!\d0_int_nxt_addr[4]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4] .extended_lut = "off";
defparam \nxt_addr[4] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[4] .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~10 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!sink0_data[60]),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[59]),
	.datae(!\int_nxt_addr_reg[4]~q ),
	.dataf(!out_data_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~10 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~10 .lut_mask = 64'h0101F1F1010FF1FF;
defparam \d0_int_nxt_addr[4]~10 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~11 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~17_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[4]~q ),
	.dataf(!\d0_int_nxt_addr[4]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~11 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~11 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[4]~11 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[1]~q ),
	.datac(!sink0_data[78]),
	.datad(!\d0_in_size[2]~1_combout ),
	.datae(!\d0_in_size[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "off";
defparam \ShiftLeft0~5 .lut_mask = 64'h000000D8000000D8;
defparam \ShiftLeft0~5 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[5] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[5]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[5] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_5),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[5]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \in_burstwrap_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[75]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[5]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[5] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[5] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[5] (
	.dataa(!new_burst_reg1),
	.datab(gnd),
	.datac(!src_payload5),
	.datad(!src_data_75),
	.datae(!\in_burstwrap_reg[5]~q ),
	.dataf(!\d0_int_nxt_addr[5]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[5] .extended_lut = "off";
defparam \nxt_addr[5] .lut_mask = 64'h00000000AAFA0050;
defparam \nxt_addr[5] .shared_arith = "off";

dffeas \int_nxt_addr_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[5]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[5] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[5]~12 (
	.dataa(!h2f_lw_ARADDR_5),
	.datab(!sink0_data[60]),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[59]),
	.datae(!\int_nxt_addr_reg[5]~q ),
	.dataf(!out_data_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[5]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[5]~12 .extended_lut = "off";
defparam \d0_int_nxt_addr[5]~12 .lut_mask = 64'h0101F1F1010FF1FF;
defparam \d0_int_nxt_addr[5]~12 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[5]~13 (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\in_burstwrap_reg[5]~q ),
	.dataf(!\d0_int_nxt_addr[5]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[5]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[5]~13 .extended_lut = "off";
defparam \d0_int_nxt_addr[5]~13 .lut_mask = 64'h00002222FFFFFFFF;
defparam \d0_int_nxt_addr[5]~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[6]~14 (
	.dataa(!h2f_lw_ARADDR_6),
	.datab(!h2f_lw_AWADDR_6),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[6]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[6]~14 .extended_lut = "off";
defparam \d0_int_nxt_addr[6]~14 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[6]~14 .shared_arith = "off";

dffeas \in_burstwrap_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[76]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[6]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[6] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[6] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[6]~8 (
	.dataa(!\int_nxt_addr_reg[6]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\in_burstwrap_reg[6]~q ),
	.datae(!\d0_int_nxt_addr[6]~14_combout ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[6]~8 .extended_lut = "off";
defparam \nxt_addr[6]~8 .lut_mask = 64'h550055000000C0C0;
defparam \nxt_addr[6]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[6]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[6]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[6] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[6] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~6 (
	.dataa(!new_burst_reg1),
	.datab(!\in_size_reg[1]~q ),
	.datac(!sink0_data[78]),
	.datad(!\d0_in_size[2]~1_combout ),
	.datae(!\d0_in_size[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~6 .extended_lut = "off";
defparam \ShiftLeft0~6 .lut_mask = 64'h0027000000270000;
defparam \ShiftLeft0~6 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[6] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[6]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[6] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_6),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[6]~q ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[6]~15 (
	.dataa(!new_burst_reg1),
	.datab(!\d0_int_nxt_addr[6]~14_combout ),
	.datac(!\int_nxt_addr_reg[6]~q ),
	.datad(!\in_burstwrap_reg[6]~q ),
	.datae(!\Add0~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[6]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[6]~15 .extended_lut = "off";
defparam \d0_int_nxt_addr[6]~15 .lut_mask = 64'h1B1B1BBB1B1B1BBB;
defparam \d0_int_nxt_addr[6]~15 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[7]~16 (
	.dataa(!h2f_lw_ARADDR_7),
	.datab(!h2f_lw_AWADDR_7),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[7]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[7]~16 .extended_lut = "off";
defparam \d0_int_nxt_addr[7]~16 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[7]~16 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[7]~7 (
	.dataa(!\int_nxt_addr_reg[7]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[7]~16_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[7]~7 .extended_lut = "off";
defparam \nxt_addr[7]~7 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[7]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg[7] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[7]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[7]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[7] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[7]~17 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[7]~16_combout ),
	.datad(!\int_nxt_addr_reg[7]~q ),
	.datae(!\Add0~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[7]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[7]~17 .extended_lut = "off";
defparam \d0_int_nxt_addr[7]~17 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[7]~17 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[8]~18 (
	.dataa(!h2f_lw_ARADDR_8),
	.datab(!h2f_lw_AWADDR_8),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[8]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[8]~18 .extended_lut = "off";
defparam \d0_int_nxt_addr[8]~18 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[8]~18 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[8]~6 (
	.dataa(!\int_nxt_addr_reg[8]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[8]~18_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[8]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[8]~6 .extended_lut = "off";
defparam \nxt_addr[8]~6 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[8]~6 .shared_arith = "off";

dffeas \int_nxt_addr_reg[8] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[8]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[8]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[8] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[8]~19 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[8]~18_combout ),
	.datad(!\int_nxt_addr_reg[8]~q ),
	.datae(!\Add0~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[8]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[8]~19 .extended_lut = "off";
defparam \d0_int_nxt_addr[8]~19 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[8]~19 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[9]~20 (
	.dataa(!h2f_lw_ARADDR_9),
	.datab(!h2f_lw_AWADDR_9),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[9]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[9]~20 .extended_lut = "off";
defparam \d0_int_nxt_addr[9]~20 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[9]~20 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[9]~5 (
	.dataa(!\int_nxt_addr_reg[9]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[9]~20_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[9]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[9]~5 .extended_lut = "off";
defparam \nxt_addr[9]~5 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[9]~5 .shared_arith = "off";

dffeas \int_nxt_addr_reg[9] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[9]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[9]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[9] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[9]~21 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[9]~20_combout ),
	.datad(!\int_nxt_addr_reg[9]~q ),
	.datae(!\Add0~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[9]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[9]~21 .extended_lut = "off";
defparam \d0_int_nxt_addr[9]~21 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[9]~21 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[10]~22 (
	.dataa(!h2f_lw_ARADDR_10),
	.datab(!h2f_lw_AWADDR_10),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[10]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[10]~22 .extended_lut = "off";
defparam \d0_int_nxt_addr[10]~22 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[10]~22 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[10]~4 (
	.dataa(!\int_nxt_addr_reg[10]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[10]~22_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[10]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[10]~4 .extended_lut = "off";
defparam \nxt_addr[10]~4 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[10]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[10] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[10]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[10]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[10] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[10]~23 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[10]~22_combout ),
	.datad(!\int_nxt_addr_reg[10]~q ),
	.datae(!\Add0~41_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[10]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[10]~23 .extended_lut = "off";
defparam \d0_int_nxt_addr[10]~23 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[10]~23 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[11]~24 (
	.dataa(!h2f_lw_ARADDR_11),
	.datab(!h2f_lw_AWADDR_11),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[11]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[11]~24 .extended_lut = "off";
defparam \d0_int_nxt_addr[11]~24 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[11]~24 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[11]~3 (
	.dataa(!\int_nxt_addr_reg[11]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[11]~24_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[11]~3 .extended_lut = "off";
defparam \nxt_addr[11]~3 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[11]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg[11] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[11]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[11]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[11] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[11] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[11]~25 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[11]~24_combout ),
	.datad(!\int_nxt_addr_reg[11]~q ),
	.datae(!\Add0~45_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[11]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[11]~25 .extended_lut = "off";
defparam \d0_int_nxt_addr[11]~25 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[11]~25 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[12]~26 (
	.dataa(!h2f_lw_ARADDR_12),
	.datab(!h2f_lw_AWADDR_12),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[12]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[12]~26 .extended_lut = "off";
defparam \d0_int_nxt_addr[12]~26 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[12]~26 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[12]~2 (
	.dataa(!\int_nxt_addr_reg[12]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[12]~26_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[12]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[12]~2 .extended_lut = "off";
defparam \nxt_addr[12]~2 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[12]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg[12] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[12]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[12]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[12] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[12] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[12]~27 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[12]~26_combout ),
	.datad(!\int_nxt_addr_reg[12]~q ),
	.datae(!\Add0~49_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[12]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[12]~27 .extended_lut = "off";
defparam \d0_int_nxt_addr[12]~27 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[12]~27 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[13]~28 (
	.dataa(!h2f_lw_ARADDR_13),
	.datab(!h2f_lw_AWADDR_13),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[13]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[13]~28 .extended_lut = "off";
defparam \d0_int_nxt_addr[13]~28 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[13]~28 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[13]~1 (
	.dataa(!\int_nxt_addr_reg[13]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[13]~28_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[13]~1 .extended_lut = "off";
defparam \nxt_addr[13]~1 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[13]~1 .shared_arith = "off";

dffeas \int_nxt_addr_reg[13] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[13]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[13]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[13] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[13] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[13]~29 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[13]~28_combout ),
	.datad(!\int_nxt_addr_reg[13]~q ),
	.datae(!\Add0~53_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[13]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[13]~29 .extended_lut = "off";
defparam \d0_int_nxt_addr[13]~29 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[13]~29 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[14]~30 (
	.dataa(!h2f_lw_ARADDR_14),
	.datab(!h2f_lw_AWADDR_14),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!sop_enable),
	.dataf(!address_burst_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[14]~30 .extended_lut = "off";
defparam \d0_int_nxt_addr[14]~30 .lut_mask = 64'h05370505053705FF;
defparam \d0_int_nxt_addr[14]~30 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[14]~0 (
	.dataa(!\int_nxt_addr_reg[14]~q ),
	.datab(!src_data_761),
	.datac(!src_data_76),
	.datad(!\d0_int_nxt_addr[14]~30_combout ),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!new_burst_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[14]~0 .extended_lut = "off";
defparam \nxt_addr[14]~0 .lut_mask = 64'h5555000000C000C0;
defparam \nxt_addr[14]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[14] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[14]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[14]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[14] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[14] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[14]~31 (
	.dataa(!new_burst_reg1),
	.datab(!\in_burstwrap_reg[6]~q ),
	.datac(!\d0_int_nxt_addr[14]~30_combout ),
	.datad(!\int_nxt_addr_reg[14]~q ),
	.datae(!\Add0~57_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[14]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[14]~31 .extended_lut = "off";
defparam \d0_int_nxt_addr[14]~31 .lut_mask = 64'h05AF27AF05AF27AF;
defparam \d0_int_nxt_addr[14]~31 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~5 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~0_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~5 .lut_mask = 64'h7777777777777777;
defparam \nxt_uncomp_subburst_byte_cnt[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~6 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~6 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~6 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~7 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~8 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~1_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~8 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~8 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~8 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~9 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~3_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~9 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~9 .lut_mask = 64'h7777777777777777;
defparam \nxt_uncomp_subburst_byte_cnt[6]~9 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_address_alignment_1 (
	ShiftLeft0,
	d0_in_size_0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	ShiftLeft0;
input 	d0_in_size_0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!ShiftLeft0),
	.datab(!d0_in_size_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4444444444444444;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_slave_agent (
	outclk_wire_0,
	mem_used_1,
	in_ready_hold,
	in_narrow_reg,
	source0_data_33,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	source0_data_35,
	in_byteen_reg_3,
	source0_data_351,
	in_byteen_reg_1,
	source0_data_331,
	WideOr0,
	out_valid_reg,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	always0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	source_endofpacket,
	in_data_reg_59,
	m0_write,
	m0_write1,
	altera_reset_synchronizer_int_chain_out,
	comb,
	WideOr01,
	cp_ready)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	mem_used_1;
input 	in_ready_hold;
input 	in_narrow_reg;
input 	source0_data_33;
input 	in_byteen_reg_2;
input 	source0_data_34;
input 	in_byteen_reg_0;
input 	source0_data_32;
input 	source0_data_35;
input 	in_byteen_reg_3;
input 	source0_data_351;
input 	in_byteen_reg_1;
input 	source0_data_331;
output 	WideOr0;
input 	out_valid_reg;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
output 	always0;
input 	mem_57_0;
input 	mem_113_0;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
output 	source_endofpacket;
input 	in_data_reg_59;
output 	m0_write;
output 	m0_write1;
input 	altera_reset_synchronizer_int_chain_out;
output 	comb;
input 	WideOr01;
output 	cp_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~0_combout ;


soc_system_altera_merlin_burst_uncompressor uncompressor(
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_used_0(mem_used_0),
	.mem_112_0(mem_112_0),
	.mem_used_01(mem_used_01),
	.always0(always0),
	.mem_57_0(mem_57_0),
	.mem_113_0(mem_113_0),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat(last_packet_beat),
	.source_endofpacket1(source_endofpacket),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(WideOr01));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!source0_data_33),
	.datab(!source0_data_32),
	.datac(!source0_data_35),
	.datad(!source0_data_351),
	.datae(!source0_data_331),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'h2222222222222222;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!source0_data_34),
	.datab(!WideOr0),
	.datac(!in_data_reg_59),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'h0007000700070007;
defparam \m0_write~1 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h8080808080808080;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!in_ready_hold),
	.datad(!\cp_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h0A8A0A8A0A8A0A8A;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_byteen_reg_1),
	.datab(!in_byteen_reg_0),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~0 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_burst_uncompressor (
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	always0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	source_endofpacket1,
	reset,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
output 	always0;
input 	mem_57_0;
input 	mem_113_0;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
output 	source_endofpacket1;
input 	reset;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~1_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \last_packet_beat~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~1_combout ;


cyclonev_lcell_comb \always0~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always0),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h007F007F007F007F;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!always0),
	.datab(!mem_57_0),
	.datac(!\burst_uncompress_busy~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!\last_packet_beat~0_combout ),
	.dataf(!\last_packet_beat~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3333333222222222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb source_endofpacket(
	.dataa(!mem_113_0),
	.datab(!last_packet_beat),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_endofpacket1),
	.sumout(),
	.cout(),
	.shareout());
defparam source_endofpacket.extended_lut = "off";
defparam source_endofpacket.lut_mask = 64'h4444444444444444;
defparam source_endofpacket.shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!always0),
	.datab(!WideOr0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'h1111111111111111;
defparam \always0~1 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~0_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_slave_translator (
	clk,
	in_ready_hold,
	source0_data_34,
	WideOr0,
	read_latency_shift_reg_0,
	m0_write,
	reset,
	in_data_reg_60)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	in_ready_hold;
input 	source0_data_34;
input 	WideOr0;
output 	read_latency_shift_reg_0;
input 	m0_write;
input 	reset;
input 	in_data_reg_60;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!in_ready_hold),
	.datab(!source0_data_34),
	.datac(!WideOr0),
	.datad(!m0_write),
	.datae(!in_data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0000001500000015;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module soc_system_soc_system_mm_interconnect_0_cmd_mux (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	Add45,
	Add55,
	Add56,
	Add46,
	nxt_out_eop,
	saved_grant_1,
	new_burst_reg,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	sink1_ready1,
	nxt_in_ready3,
	saved_grant_0,
	src_valid,
	altera_reset_synchronizer_int_chain_out,
	WideOr11,
	src_payload_0,
	src_data_78,
	src_data_79,
	src_data_77,
	src_payload,
	Add1,
	log2ceil,
	src_payload1,
	Add3,
	log2ceil1,
	src_data_71,
	src_payload2,
	log2ceil2,
	src_payload3,
	Add31,
	src_data_70,
	src_data_34,
	src_data_32,
	src_data_35,
	src_data_33,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_72,
	src_payload7,
	Selector17,
	src_data_73,
	src_payload8,
	src_payload9,
	src_data_74,
	src_payload10,
	src_payload11,
	src_data_75,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_data_711,
	src_data_701,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_721,
	src_data_731,
	src_data_741,
	src_data_751,
	src_data_76,
	src_data_761,
	src_data_762)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	Add4;
input 	Add5;
input 	Add41;
input 	Add51;
input 	Add42;
input 	Add52;
input 	Add43;
input 	Add53;
input 	Add44;
input 	Add54;
input 	Add45;
input 	Add55;
input 	Add56;
input 	Add46;
input 	nxt_out_eop;
output 	saved_grant_1;
input 	new_burst_reg;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
output 	sink1_ready1;
input 	nxt_in_ready3;
output 	saved_grant_0;
output 	src_valid;
input 	altera_reset_synchronizer_int_chain_out;
output 	WideOr11;
output 	src_payload_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_77;
output 	src_payload;
input 	Add1;
input 	log2ceil;
output 	src_payload1;
input 	Add3;
input 	log2ceil1;
output 	src_data_71;
output 	src_payload2;
input 	log2ceil2;
output 	src_payload3;
input 	Add31;
output 	src_data_70;
output 	src_data_34;
output 	src_data_32;
output 	src_data_35;
output 	src_data_33;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_data_72;
output 	src_payload7;
input 	Selector17;
output 	src_data_73;
output 	src_payload8;
output 	src_payload9;
output 	src_data_74;
output 	src_payload10;
output 	src_payload11;
output 	src_data_75;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_data_711;
output 	src_data_701;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_721;
output 	src_data_731;
output 	src_data_741;
output 	src_data_751;
output 	src_data_76;
output 	src_data_761;
output 	src_data_762;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_payload~1_combout ;
wire \src_payload~3_combout ;
wire \src_data[73]~0_combout ;
wire \src_data[71]~1_combout ;
wire \src_data[70]~2_combout ;
wire \src_data[74]~4_combout ;
wire \src_data[70]~5_combout ;
wire \src_data[72]~7_combout ;
wire \src_data[72]~8_combout ;
wire \src_data[73]~10_combout ;
wire \src_data[74]~12_combout ;
wire \src_data[75]~14_combout ;
wire \src_data[76]~24_combout ;


soc_system_altera_merlin_arbitrator arb(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.clk(outclk_wire_0),
	.nxt_in_ready(nxt_in_ready3),
	.grant_1(\arb|grant[1]~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr1(WideOr11),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ));

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb sink1_ready(
	.dataa(!saved_grant_1),
	.datab(!new_burst_reg),
	.datac(!nxt_in_ready),
	.datad(!nxt_out_eop),
	.datae(!nxt_in_ready1),
	.dataf(!nxt_in_ready2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink1_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam sink1_ready.extended_lut = "off";
defparam sink1_ready.lut_mask = 64'h0105555555555555;
defparam sink1_ready.shared_arith = "off";

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0101010101010101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!saved_grant_1),
	.datae(!saved_grant_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0055035700550357;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h0202020202020202;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!Add1),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h8000000080000000;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~3 (
	.dataa(!Add5),
	.datab(!\src_payload~1_combout ),
	.datac(!src_payload1),
	.datad(!\src_payload~3_combout ),
	.datae(!\src_data[71]~1_combout ),
	.dataf(!\src_data[70]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~3 .extended_lut = "off";
defparam \src_data[71]~3 .lut_mask = 64'hEE0E000000000000;
defparam \src_data[71]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add41),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h0202020202020202;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!h2f_lw_AWSIZE_1),
	.datad(!h2f_lw_AWSIZE_2),
	.datae(!log2ceil2),
	.dataf(!log2ceil),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h8000000000000000;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~6 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~3_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add51),
	.datae(!src_payload3),
	.dataf(!\src_data[70]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~6 .extended_lut = "off";
defparam \src_data[70]~6 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[70]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add42),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h0202020202020202;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!h2f_lw_AWSIZE_1),
	.datad(!h2f_lw_AWSIZE_2),
	.datae(!log2ceil2),
	.dataf(!log2ceil),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'hA800A00080000000;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~9 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~3_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add52),
	.datae(!src_payload6),
	.dataf(!\src_data[72]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~9 .extended_lut = "off";
defparam \src_data[72]~9 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[72]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add43),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h0202020202020202;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~11 (
	.dataa(!\src_payload~1_combout ),
	.datab(!Selector17),
	.datac(!\src_payload~3_combout ),
	.datad(!Add53),
	.datae(!\src_data[73]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~11 .extended_lut = "off";
defparam \src_data[73]~11 .lut_mask = 64'h0000F3A20000F3A2;
defparam \src_data[73]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add44),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0202020202020202;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!h2f_lw_AWSIZE_1),
	.datad(!h2f_lw_AWSIZE_2),
	.datae(!log2ceil2),
	.dataf(!log2ceil),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'hEA80AA00A800A000;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~13 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~3_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add54),
	.datae(!src_payload9),
	.dataf(!\src_data[74]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~13 .extended_lut = "off";
defparam \src_data[74]~13 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[74]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(!Add45),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h0202020202020202;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!Add1),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'hE8A0A080E8A0A080;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[75]~15 (
	.dataa(!\src_payload~1_combout ),
	.datab(!\src_payload~3_combout ),
	.datac(!\src_data[70]~2_combout ),
	.datad(!Add55),
	.datae(!src_payload11),
	.dataf(!\src_data[75]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_75),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[75]~15 .extended_lut = "off";
defparam \src_data[75]~15 .lut_mask = 64'hC080F0A000000000;
defparam \src_data[75]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h1111111111111111;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h1111111111111111;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'h1111111111111111;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'h1111111111111111;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~36 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~36 .extended_lut = "off";
defparam \src_payload~36 .lut_mask = 64'h1111111111111111;
defparam \src_payload~36 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~37 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~37 .extended_lut = "off";
defparam \src_payload~37 .lut_mask = 64'h1111111111111111;
defparam \src_payload~37 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~38 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload36),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~38 .extended_lut = "off";
defparam \src_payload~38 .lut_mask = 64'h1111111111111111;
defparam \src_payload~38 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~39 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload37),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~39 .extended_lut = "off";
defparam \src_payload~39 .lut_mask = 64'h1111111111111111;
defparam \src_payload~39 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~40 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~40 .extended_lut = "off";
defparam \src_payload~40 .lut_mask = 64'h1111111111111111;
defparam \src_payload~40 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~41 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~41 .extended_lut = "off";
defparam \src_payload~41 .lut_mask = 64'h1111111111111111;
defparam \src_payload~41 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~42 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~42 .extended_lut = "off";
defparam \src_payload~42 .lut_mask = 64'h1111111111111111;
defparam \src_payload~42 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~43 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~43 .extended_lut = "off";
defparam \src_payload~43 .lut_mask = 64'h1111111111111111;
defparam \src_payload~43 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~44 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~44 .extended_lut = "off";
defparam \src_payload~44 .lut_mask = 64'h1111111111111111;
defparam \src_payload~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~16 (
	.dataa(!src_payload),
	.datab(!src_data_71),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_711),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~16 .extended_lut = "off";
defparam \src_data[71]~16 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[71]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~17 (
	.dataa(!src_payload2),
	.datab(!src_data_70),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_701),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~17 .extended_lut = "off";
defparam \src_data[70]~17 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[70]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~18 (
	.dataa(!src_payload5),
	.datab(!src_data_72),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_721),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~18 .extended_lut = "off";
defparam \src_data[72]~18 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[72]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~19 (
	.dataa(!src_payload7),
	.datab(!src_data_73),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_731),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~19 .extended_lut = "off";
defparam \src_data[73]~19 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[73]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~20 (
	.dataa(!src_payload8),
	.datab(!src_data_74),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_741),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~20 .extended_lut = "off";
defparam \src_data[74]~20 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[74]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[75]~21 (
	.dataa(!src_payload10),
	.datab(!src_data_75),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_751),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[75]~21 .extended_lut = "off";
defparam \src_data[75]~21 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \src_data[75]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~22 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add56),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_76),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~22 .extended_lut = "off";
defparam \src_data[76]~22 .lut_mask = 64'h050D050D050D050D;
defparam \src_data[76]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~23 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!Add46),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_761),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~23 .extended_lut = "off";
defparam \src_data[76]~23 .lut_mask = 64'h050D050D050D050D;
defparam \src_data[76]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~25 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!Add56),
	.dataf(!\src_data[76]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_762),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~25 .extended_lut = "off";
defparam \src_data[76]~25 .lut_mask = 64'h05FF0DFF05050D0D;
defparam \src_data[76]~25 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready3),
	.datab(!WideOr11),
	.datac(!src_payload_0),
	.datad(!\packet_in_progress~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hCE02CE02CE02CE02;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h2222222222222222;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_AWBURST_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~0 (
	.dataa(!h2f_lw_ARBURST_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~0 .extended_lut = "off";
defparam \src_data[73]~0 .lut_mask = 64'h1111111111111111;
defparam \src_data[73]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~1 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!\src_data[73]~0_combout ),
	.datae(!Add3),
	.dataf(!log2ceil1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~1 .extended_lut = "off";
defparam \src_data[71]~1 .lut_mask = 64'h00FF00FF007F00FF;
defparam \src_data[71]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~2 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_AWBURST_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~2 .extended_lut = "off";
defparam \src_data[70]~2 .lut_mask = 64'h0537053705370537;
defparam \src_data[70]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~4 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~4 .extended_lut = "off";
defparam \src_data[74]~4 .lut_mask = 64'h80FF0F0030004000;
defparam \src_data[74]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~5 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\src_data[73]~0_combout ),
	.datad(!Add31),
	.datae(!\src_data[74]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~5 .extended_lut = "off";
defparam \src_data[70]~5 .lut_mask = 64'h0F0F070F0F0F070F;
defparam \src_data[70]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~7 .extended_lut = "off";
defparam \src_data[72]~7 .lut_mask = 64'h0F003000400080FF;
defparam \src_data[72]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~8 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\src_data[73]~0_combout ),
	.datad(!Add31),
	.datae(!\src_data[72]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~8 .extended_lut = "off";
defparam \src_data[72]~8 .lut_mask = 64'h070F0F0F070F0F0F;
defparam \src_data[72]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~10 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\src_data[73]~0_combout ),
	.datad(!Add31),
	.datae(!\src_data[70]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~10 .extended_lut = "off";
defparam \src_data[73]~10 .lut_mask = 64'hF8F00000F8F00000;
defparam \src_data[73]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~12 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\src_data[73]~0_combout ),
	.datad(!Add31),
	.datae(!\src_data[74]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~12 .extended_lut = "off";
defparam \src_data[74]~12 .lut_mask = 64'h070F0107070F0107;
defparam \src_data[74]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[75]~14 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(!\src_data[73]~0_combout ),
	.datae(!Add3),
	.dataf(!log2ceil1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[75]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[75]~14 .extended_lut = "off";
defparam \src_data[75]~14 .lut_mask = 64'h001F007F0017005F;
defparam \src_data[75]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~24 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Add46),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[76]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~24 .extended_lut = "off";
defparam \src_data[76]~24 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \src_data[76]~24 .shared_arith = "off";

endmodule

module soc_system_altera_merlin_arbitrator (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	clk,
	nxt_in_ready,
	grant_1,
	reset,
	WideOr1,
	src_payload_0,
	packet_in_progress,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	clk;
input 	nxt_in_ready;
output 	grant_1;
input 	reset;
input 	WideOr1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h5455005554550055;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0303000203030002;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hA8A8A8A8A8A8A8A8;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready),
	.datab(!WideOr1),
	.datac(!src_payload_0),
	.datad(!packet_in_progress),
	.datae(!\top_priority_reg[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hCE020000CE020000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module soc_system_soc_system_mm_interconnect_0_rsp_demux (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	always0,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src0_valid2,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	always0;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src0_valid2;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_59_0),
	.datab(!mem_57_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!always0),
	.datad(!src0_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h007F007F007F007F;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!always0),
	.datad(!src0_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F007F007F007F00;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!src0_valid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3535353535353535;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module soc_system_soc_system_onchip_memory2_0 (
	outclk_wire_0,
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	q_a_16,
	q_b_16,
	q_a_17,
	q_b_17,
	q_a_18,
	q_b_18,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	q_a_21,
	q_b_21,
	q_a_22,
	q_b_22,
	q_a_23,
	q_b_23,
	q_a_24,
	q_b_24,
	q_a_25,
	q_b_25,
	q_a_26,
	q_b_26,
	q_a_27,
	q_b_27,
	q_a_28,
	q_b_28,
	q_a_29,
	q_b_29,
	q_a_30,
	q_b_30,
	q_a_31,
	q_b_31,
	source0_data_34,
	source0_data_32,
	m0_write,
	in_data_reg_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	int_nxt_addr_reg_dly_10,
	int_nxt_addr_reg_dly_11,
	int_nxt_addr_reg_dly_12,
	int_nxt_addr_reg_dly_13,
	int_nxt_addr_reg_dly_14,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	source0_data_33,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	source0_data_35,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	ram_mm_chipselect,
	ram_mm_write,
	ram_clk_clk,
	ram_mm_clken,
	ram_mm_writedata_0,
	ram_mm_address_0,
	ram_mm_address_1,
	ram_mm_address_2,
	ram_mm_address_3,
	ram_mm_address_4,
	ram_mm_address_5,
	ram_mm_address_6,
	ram_mm_address_7,
	ram_mm_address_8,
	ram_mm_address_9,
	ram_mm_address_10,
	ram_mm_address_11,
	ram_mm_address_12,
	ram_mm_byteenable_0,
	ram_mm_writedata_1,
	ram_mm_writedata_2,
	ram_mm_writedata_3,
	ram_mm_writedata_4,
	ram_mm_writedata_5,
	ram_mm_writedata_6,
	ram_mm_writedata_7,
	ram_mm_writedata_8,
	ram_mm_byteenable_1,
	ram_mm_writedata_9,
	ram_mm_writedata_10,
	ram_mm_writedata_11,
	ram_mm_writedata_12,
	ram_mm_writedata_13,
	ram_mm_writedata_14,
	ram_mm_writedata_15,
	ram_mm_writedata_16,
	ram_mm_byteenable_2,
	ram_mm_writedata_17,
	ram_mm_writedata_18,
	ram_mm_writedata_19,
	ram_mm_writedata_20,
	ram_mm_writedata_21,
	ram_mm_writedata_22,
	ram_mm_writedata_23,
	ram_mm_writedata_24,
	ram_mm_byteenable_3,
	ram_mm_writedata_25,
	ram_mm_writedata_26,
	ram_mm_writedata_27,
	ram_mm_writedata_28,
	ram_mm_writedata_29,
	ram_mm_writedata_30,
	ram_mm_writedata_31)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
output 	q_a_8;
output 	q_b_8;
output 	q_a_9;
output 	q_b_9;
output 	q_a_10;
output 	q_b_10;
output 	q_a_11;
output 	q_b_11;
output 	q_a_12;
output 	q_b_12;
output 	q_a_13;
output 	q_b_13;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
output 	q_a_16;
output 	q_b_16;
output 	q_a_17;
output 	q_b_17;
output 	q_a_18;
output 	q_b_18;
output 	q_a_19;
output 	q_b_19;
output 	q_a_20;
output 	q_b_20;
output 	q_a_21;
output 	q_b_21;
output 	q_a_22;
output 	q_b_22;
output 	q_a_23;
output 	q_b_23;
output 	q_a_24;
output 	q_b_24;
output 	q_a_25;
output 	q_b_25;
output 	q_a_26;
output 	q_b_26;
output 	q_a_27;
output 	q_b_27;
output 	q_a_28;
output 	q_b_28;
output 	q_a_29;
output 	q_b_29;
output 	q_a_30;
output 	q_b_30;
output 	q_a_31;
output 	q_b_31;
input 	source0_data_34;
input 	source0_data_32;
input 	m0_write;
input 	in_data_reg_0;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_5;
input 	int_nxt_addr_reg_dly_6;
input 	int_nxt_addr_reg_dly_7;
input 	int_nxt_addr_reg_dly_8;
input 	int_nxt_addr_reg_dly_9;
input 	int_nxt_addr_reg_dly_10;
input 	int_nxt_addr_reg_dly_11;
input 	int_nxt_addr_reg_dly_12;
input 	int_nxt_addr_reg_dly_13;
input 	int_nxt_addr_reg_dly_14;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	source0_data_33;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	source0_data_35;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
input 	ram_mm_chipselect;
input 	ram_mm_write;
input 	ram_clk_clk;
input 	ram_mm_clken;
input 	ram_mm_writedata_0;
input 	ram_mm_address_0;
input 	ram_mm_address_1;
input 	ram_mm_address_2;
input 	ram_mm_address_3;
input 	ram_mm_address_4;
input 	ram_mm_address_5;
input 	ram_mm_address_6;
input 	ram_mm_address_7;
input 	ram_mm_address_8;
input 	ram_mm_address_9;
input 	ram_mm_address_10;
input 	ram_mm_address_11;
input 	ram_mm_address_12;
input 	ram_mm_byteenable_0;
input 	ram_mm_writedata_1;
input 	ram_mm_writedata_2;
input 	ram_mm_writedata_3;
input 	ram_mm_writedata_4;
input 	ram_mm_writedata_5;
input 	ram_mm_writedata_6;
input 	ram_mm_writedata_7;
input 	ram_mm_writedata_8;
input 	ram_mm_byteenable_1;
input 	ram_mm_writedata_9;
input 	ram_mm_writedata_10;
input 	ram_mm_writedata_11;
input 	ram_mm_writedata_12;
input 	ram_mm_writedata_13;
input 	ram_mm_writedata_14;
input 	ram_mm_writedata_15;
input 	ram_mm_writedata_16;
input 	ram_mm_byteenable_2;
input 	ram_mm_writedata_17;
input 	ram_mm_writedata_18;
input 	ram_mm_writedata_19;
input 	ram_mm_writedata_20;
input 	ram_mm_writedata_21;
input 	ram_mm_writedata_22;
input 	ram_mm_writedata_23;
input 	ram_mm_writedata_24;
input 	ram_mm_byteenable_3;
input 	ram_mm_writedata_25;
input 	ram_mm_writedata_26;
input 	ram_mm_writedata_27;
input 	ram_mm_writedata_28;
input 	ram_mm_writedata_29;
input 	ram_mm_writedata_30;
input 	ram_mm_writedata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren2~combout ;


soc_system_altsyncram_1 the_altsyncram(
	.clock0(outclk_wire_0),
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.byteena_a({source0_data_35,source0_data_34,source0_data_33,source0_data_32}),
	.wren_a(m0_write),
	.wren_b(\wren2~combout ),
	.data_a({in_data_reg_31,in_data_reg_30,in_data_reg_29,in_data_reg_28,in_data_reg_27,in_data_reg_26,in_data_reg_25,in_data_reg_24,in_data_reg_23,in_data_reg_22,in_data_reg_21,in_data_reg_20,in_data_reg_19,in_data_reg_18,in_data_reg_17,in_data_reg_16,in_data_reg_15,in_data_reg_14,
in_data_reg_13,in_data_reg_12,in_data_reg_11,in_data_reg_10,in_data_reg_9,in_data_reg_8,in_data_reg_7,in_data_reg_6,in_data_reg_5,in_data_reg_4,in_data_reg_3,in_data_reg_2,in_data_reg_1,in_data_reg_0}),
	.address_a({int_nxt_addr_reg_dly_14,int_nxt_addr_reg_dly_13,int_nxt_addr_reg_dly_12,int_nxt_addr_reg_dly_11,int_nxt_addr_reg_dly_10,int_nxt_addr_reg_dly_9,int_nxt_addr_reg_dly_8,int_nxt_addr_reg_dly_7,int_nxt_addr_reg_dly_6,int_nxt_addr_reg_dly_5,int_nxt_addr_reg_dly_4,
int_nxt_addr_reg_dly_3,int_nxt_addr_reg_dly_2}),
	.clock1(ram_clk_clk),
	.clocken1(ram_mm_clken),
	.data_b({ram_mm_writedata_31,ram_mm_writedata_30,ram_mm_writedata_29,ram_mm_writedata_28,ram_mm_writedata_27,ram_mm_writedata_26,ram_mm_writedata_25,ram_mm_writedata_24,ram_mm_writedata_23,ram_mm_writedata_22,ram_mm_writedata_21,ram_mm_writedata_20,ram_mm_writedata_19,
ram_mm_writedata_18,ram_mm_writedata_17,ram_mm_writedata_16,ram_mm_writedata_15,ram_mm_writedata_14,ram_mm_writedata_13,ram_mm_writedata_12,ram_mm_writedata_11,ram_mm_writedata_10,ram_mm_writedata_9,ram_mm_writedata_8,ram_mm_writedata_7,ram_mm_writedata_6,
ram_mm_writedata_5,ram_mm_writedata_4,ram_mm_writedata_3,ram_mm_writedata_2,ram_mm_writedata_1,ram_mm_writedata_0}),
	.address_b({ram_mm_address_12,ram_mm_address_11,ram_mm_address_10,ram_mm_address_9,ram_mm_address_8,ram_mm_address_7,ram_mm_address_6,ram_mm_address_5,ram_mm_address_4,ram_mm_address_3,ram_mm_address_2,ram_mm_address_1,ram_mm_address_0}),
	.byteena_b({ram_mm_byteenable_3,ram_mm_byteenable_2,ram_mm_byteenable_1,ram_mm_byteenable_0}));

cyclonev_lcell_comb wren2(
	.dataa(!ram_mm_chipselect),
	.datab(!ram_mm_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren2~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wren2.extended_lut = "off";
defparam wren2.lut_mask = 64'h1111111111111111;
defparam wren2.shared_arith = "off";

endmodule

module soc_system_altsyncram_1 (
	clock0,
	q_a,
	q_b,
	byteena_a,
	wren_a,
	wren_b,
	data_a,
	address_a,
	clock1,
	clocken1,
	data_b,
	address_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	[3:0] byteena_a;
input 	wren_a;
input 	wren_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	clock1;
input 	clocken1;
input 	[31:0] data_b;
input 	[12:0] address_b;
input 	[3:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altsyncram_jcd2 auto_generated(
	.clock0(clock0),
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.wren_a(wren_a),
	.wren_b(wren_b),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock1(clock1),
	.clocken1(clocken1),
	.data_b({data_b[31],data_b[30],data_b[29],data_b[28],data_b[27],data_b[26],data_b[25],data_b[24],data_b[23],data_b[22],data_b[21],data_b[20],data_b[19],data_b[18],data_b[17],data_b[16],data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.address_b({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.byteena_b({byteena_b[3],byteena_b[2],byteena_b[1],byteena_b[0]}));

endmodule

module soc_system_altsyncram_jcd2 (
	clock0,
	q_a,
	q_b,
	byteena_a,
	wren_a,
	wren_b,
	data_a,
	address_a,
	clock1,
	clocken1,
	data_b,
	address_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	[3:0] byteena_a;
input 	wren_a;
input 	wren_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	clock1;
input 	clocken1;
input 	[31:0] data_b;
input 	[12:0] address_b;
input 	[3:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 8192;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 13;
defparam ram_block1a0.port_b_byte_enable_clock = "clock1";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock1";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 8191;
defparam ram_block1a0.port_b_logical_ram_depth = 8192;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.port_b_write_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 8192;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 13;
defparam ram_block1a1.port_b_byte_enable_clock = "clock1";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock1";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 8191;
defparam ram_block1a1.port_b_logical_ram_depth = 8192;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.port_b_write_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 8192;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 13;
defparam ram_block1a2.port_b_byte_enable_clock = "clock1";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock1";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 8191;
defparam ram_block1a2.port_b_logical_ram_depth = 8192;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.port_b_write_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 8192;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 13;
defparam ram_block1a3.port_b_byte_enable_clock = "clock1";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock1";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 8191;
defparam ram_block1a3.port_b_logical_ram_depth = 8192;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.port_b_write_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 8192;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 13;
defparam ram_block1a4.port_b_byte_enable_clock = "clock1";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock1";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 8191;
defparam ram_block1a4.port_b_logical_ram_depth = 8192;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.port_b_write_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 8192;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 13;
defparam ram_block1a5.port_b_byte_enable_clock = "clock1";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock1";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 8191;
defparam ram_block1a5.port_b_logical_ram_depth = 8192;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.port_b_write_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 8192;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 13;
defparam ram_block1a6.port_b_byte_enable_clock = "clock1";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock1";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 8191;
defparam ram_block1a6.port_b_logical_ram_depth = 8192;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.port_b_write_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 8192;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 13;
defparam ram_block1a7.port_b_byte_enable_clock = "clock1";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock1";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 8191;
defparam ram_block1a7.port_b_logical_ram_depth = 8192;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.port_b_write_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 8192;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 13;
defparam ram_block1a8.port_b_byte_enable_clock = "clock1";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock1";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 8191;
defparam ram_block1a8.port_b_logical_ram_depth = 8192;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.port_b_write_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 8192;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 13;
defparam ram_block1a9.port_b_byte_enable_clock = "clock1";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock1";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 8191;
defparam ram_block1a9.port_b_logical_ram_depth = 8192;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.port_b_write_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 8192;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 13;
defparam ram_block1a10.port_b_byte_enable_clock = "clock1";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock1";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 8191;
defparam ram_block1a10.port_b_logical_ram_depth = 8192;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.port_b_write_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 8192;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 13;
defparam ram_block1a11.port_b_byte_enable_clock = "clock1";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock1";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 8191;
defparam ram_block1a11.port_b_logical_ram_depth = 8192;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.port_b_write_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 8192;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 13;
defparam ram_block1a12.port_b_byte_enable_clock = "clock1";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock1";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 8191;
defparam ram_block1a12.port_b_logical_ram_depth = 8192;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.port_b_write_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 8192;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 13;
defparam ram_block1a13.port_b_byte_enable_clock = "clock1";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock1";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 8191;
defparam ram_block1a13.port_b_logical_ram_depth = 8192;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.port_b_write_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 8192;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 13;
defparam ram_block1a14.port_b_byte_enable_clock = "clock1";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock1";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 8191;
defparam ram_block1a14.port_b_logical_ram_depth = 8192;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.port_b_write_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 8192;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 13;
defparam ram_block1a15.port_b_byte_enable_clock = "clock1";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock1";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 8191;
defparam ram_block1a15.port_b_logical_ram_depth = 8192;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.port_b_write_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 8192;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 13;
defparam ram_block1a16.port_b_byte_enable_clock = "clock1";
defparam ram_block1a16.port_b_byte_enable_mask_width = 1;
defparam ram_block1a16.port_b_byte_size = 1;
defparam ram_block1a16.port_b_data_in_clock = "clock1";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 8191;
defparam ram_block1a16.port_b_logical_ram_depth = 8192;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.port_b_write_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 8192;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 13;
defparam ram_block1a17.port_b_byte_enable_clock = "clock1";
defparam ram_block1a17.port_b_byte_enable_mask_width = 1;
defparam ram_block1a17.port_b_byte_size = 1;
defparam ram_block1a17.port_b_data_in_clock = "clock1";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 8191;
defparam ram_block1a17.port_b_logical_ram_depth = 8192;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.port_b_write_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 8192;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 13;
defparam ram_block1a18.port_b_byte_enable_clock = "clock1";
defparam ram_block1a18.port_b_byte_enable_mask_width = 1;
defparam ram_block1a18.port_b_byte_size = 1;
defparam ram_block1a18.port_b_data_in_clock = "clock1";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 8191;
defparam ram_block1a18.port_b_logical_ram_depth = 8192;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.port_b_write_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 8192;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 13;
defparam ram_block1a19.port_b_byte_enable_clock = "clock1";
defparam ram_block1a19.port_b_byte_enable_mask_width = 1;
defparam ram_block1a19.port_b_byte_size = 1;
defparam ram_block1a19.port_b_data_in_clock = "clock1";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 8191;
defparam ram_block1a19.port_b_logical_ram_depth = 8192;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.port_b_write_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 8192;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 13;
defparam ram_block1a20.port_b_byte_enable_clock = "clock1";
defparam ram_block1a20.port_b_byte_enable_mask_width = 1;
defparam ram_block1a20.port_b_byte_size = 1;
defparam ram_block1a20.port_b_data_in_clock = "clock1";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 8191;
defparam ram_block1a20.port_b_logical_ram_depth = 8192;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.port_b_write_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 8192;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 13;
defparam ram_block1a21.port_b_byte_enable_clock = "clock1";
defparam ram_block1a21.port_b_byte_enable_mask_width = 1;
defparam ram_block1a21.port_b_byte_size = 1;
defparam ram_block1a21.port_b_data_in_clock = "clock1";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 8191;
defparam ram_block1a21.port_b_logical_ram_depth = 8192;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.port_b_write_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 8192;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 13;
defparam ram_block1a22.port_b_byte_enable_clock = "clock1";
defparam ram_block1a22.port_b_byte_enable_mask_width = 1;
defparam ram_block1a22.port_b_byte_size = 1;
defparam ram_block1a22.port_b_data_in_clock = "clock1";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 8191;
defparam ram_block1a22.port_b_logical_ram_depth = 8192;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.port_b_write_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 8192;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 13;
defparam ram_block1a23.port_b_byte_enable_clock = "clock1";
defparam ram_block1a23.port_b_byte_enable_mask_width = 1;
defparam ram_block1a23.port_b_byte_size = 1;
defparam ram_block1a23.port_b_data_in_clock = "clock1";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 8191;
defparam ram_block1a23.port_b_logical_ram_depth = 8192;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.port_b_write_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "bidir_dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 8192;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 13;
defparam ram_block1a24.port_b_byte_enable_clock = "clock1";
defparam ram_block1a24.port_b_byte_enable_mask_width = 1;
defparam ram_block1a24.port_b_byte_size = 1;
defparam ram_block1a24.port_b_data_in_clock = "clock1";
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 8191;
defparam ram_block1a24.port_b_logical_ram_depth = 8192;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.port_b_write_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "bidir_dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 8192;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 13;
defparam ram_block1a25.port_b_byte_enable_clock = "clock1";
defparam ram_block1a25.port_b_byte_enable_mask_width = 1;
defparam ram_block1a25.port_b_byte_size = 1;
defparam ram_block1a25.port_b_data_in_clock = "clock1";
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 8191;
defparam ram_block1a25.port_b_logical_ram_depth = 8192;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.port_b_write_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "bidir_dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 8192;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 13;
defparam ram_block1a26.port_b_byte_enable_clock = "clock1";
defparam ram_block1a26.port_b_byte_enable_mask_width = 1;
defparam ram_block1a26.port_b_byte_size = 1;
defparam ram_block1a26.port_b_data_in_clock = "clock1";
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 8191;
defparam ram_block1a26.port_b_logical_ram_depth = 8192;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.port_b_write_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "bidir_dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 8192;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 13;
defparam ram_block1a27.port_b_byte_enable_clock = "clock1";
defparam ram_block1a27.port_b_byte_enable_mask_width = 1;
defparam ram_block1a27.port_b_byte_size = 1;
defparam ram_block1a27.port_b_data_in_clock = "clock1";
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 8191;
defparam ram_block1a27.port_b_logical_ram_depth = 8192;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.port_b_write_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "bidir_dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 8192;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 13;
defparam ram_block1a28.port_b_byte_enable_clock = "clock1";
defparam ram_block1a28.port_b_byte_enable_mask_width = 1;
defparam ram_block1a28.port_b_byte_size = 1;
defparam ram_block1a28.port_b_data_in_clock = "clock1";
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 8191;
defparam ram_block1a28.port_b_logical_ram_depth = 8192;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.port_b_write_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "bidir_dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 8192;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 13;
defparam ram_block1a29.port_b_byte_enable_clock = "clock1";
defparam ram_block1a29.port_b_byte_enable_mask_width = 1;
defparam ram_block1a29.port_b_byte_size = 1;
defparam ram_block1a29.port_b_data_in_clock = "clock1";
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 8191;
defparam ram_block1a29.port_b_logical_ram_depth = 8192;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.port_b_write_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "bidir_dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 8192;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 13;
defparam ram_block1a30.port_b_byte_enable_clock = "clock1";
defparam ram_block1a30.port_b_byte_enable_mask_width = 1;
defparam ram_block1a30.port_b_byte_size = 1;
defparam ram_block1a30.port_b_data_in_clock = "clock1";
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 8191;
defparam ram_block1a30.port_b_logical_ram_depth = 8192;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.port_b_write_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "/home/imants/programs/git/VGA_Ambilight/soc_project/ram_memory.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "soc_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_jcd2:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "bidir_dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 8192;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 13;
defparam ram_block1a31.port_b_byte_enable_clock = "clock1";
defparam ram_block1a31.port_b_byte_enable_mask_width = 1;
defparam ram_block1a31.port_b_byte_size = 1;
defparam ram_block1a31.port_b_data_in_clock = "clock1";
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 8191;
defparam ram_block1a31.port_b_logical_ram_depth = 8192;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.port_b_write_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

endmodule

module soc_system_soc_system_pll_0 (
	outclk_wire_0,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_0;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



soc_system_altera_pll_1 altera_pll_i(
	.outclk({outclk_wire_0}),
	.refclk(clk_clk),
	.rst(reset_reset_n));

endmodule

module soc_system_altera_pll_1 (
	outclk,
	refclk,
	rst)/* synthesis synthesis_greybox=0 */;
output 	[0:0] outclk;
input 	refclk;
input 	rst;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fboutclk_wire[0] ;


generic_pll \general[0].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(!rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[0]),
	.fboutclk(\fboutclk_wire[0] ),
	.locked(),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[0].gpll .clock_name_global = "false";
defparam \general[0].gpll .duty_cycle = 50;
defparam \general[0].gpll .fractional_vco_multiplier = "false";
defparam \general[0].gpll .output_clock_frequency = "100.0 mhz";
defparam \general[0].gpll .phase_shift = "0 ps";
defparam \general[0].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[0].gpll .simulation_type = "timing";

endmodule
