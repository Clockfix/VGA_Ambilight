ram2port_inst : ram2port PORT MAP(
	clock => clock_sig,
	data => data_sig,
	rdaddress => rdaddress_sig,
	rden => rden_sig,
	wraddress => wraddress_sig,
	wren => wren_sig,
	q => q_sig
);